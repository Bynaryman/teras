* NGSPICE file created from teras.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

.subckt teras VGND VPWR clk data_i[0] data_i[10] data_i[11] data_i[12] data_i[13]
+ data_i[14] data_i[15] data_i[16] data_i[17] data_i[18] data_i[19] data_i[1] data_i[20]
+ data_i[21] data_i[22] data_i[23] data_i[24] data_i[25] data_i[26] data_i[27] data_i[28]
+ data_i[29] data_i[2] data_i[30] data_i[31] data_i[3] data_i[4] data_i[5] data_i[6]
+ data_i[7] data_i[8] data_i[9] data_o[0] data_o[10] data_o[11] data_o[12] data_o[13]
+ data_o[14] data_o[15] data_o[16] data_o[17] data_o[18] data_o[19] data_o[1] data_o[20]
+ data_o[21] data_o[22] data_o[23] data_o[24] data_o[25] data_o[26] data_o[27] data_o[28]
+ data_o[29] data_o[2] data_o[30] data_o[31] data_o[3] data_o[4] data_o[5] data_o[6]
+ data_o[7] data_o[8] data_o[9] rst_n rtr_i rtr_o rts_i rts_o
XFILLER_67_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05903_ _05903_/A _05903_/B _05903_/C VGND VGND VPWR VPWR _05904_/D sky130_fd_sc_hd__or3_1
XFILLER_28_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06883_ _07962_/B VGND VGND VPWR VPWR _07955_/B sky130_fd_sc_hd__clkbuf_2
X_09671_ _09671_/A _09671_/B VGND VGND VPWR VPWR _13667_/D sky130_fd_sc_hd__xor2_1
XFILLER_67_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08622_ _08622_/A _08622_/B VGND VGND VPWR VPWR _08622_/X sky130_fd_sc_hd__or2_1
XFILLER_54_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08553_ _08567_/A _08582_/B VGND VGND VPWR VPWR _09407_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07504_ _07504_/A _07504_/B _07504_/C _07504_/D VGND VGND VPWR VPWR _07533_/A sky130_fd_sc_hd__or4_1
X_08484_ _08733_/A VGND VGND VPWR VPWR _08642_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_35_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07435_ _07435_/A _07435_/B VGND VGND VPWR VPWR _09177_/B sky130_fd_sc_hd__nand2_1
XFILLER_149_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07366_ _13139_/Q _09130_/B VGND VGND VPWR VPWR _07416_/A sky130_fd_sc_hd__xnor2_1
XFILLER_149_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06317_ hold199/A _14184_/D _14185_/D _14188_/D VGND VGND VPWR VPWR _06318_/D sky130_fd_sc_hd__or4_1
X_09105_ _09105_/A VGND VGND VPWR VPWR _13526_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07297_ _07297_/A VGND VGND VPWR VPWR _13134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09036_ _13218_/Q _13447_/Q _09040_/S VGND VGND VPWR VPWR _09037_/A sky130_fd_sc_hd__mux2_1
X_06248_ _06248_/A VGND VGND VPWR VPWR _14393_/D sky130_fd_sc_hd__clkbuf_1
Xhold340 hold340/A VGND VGND VPWR VPWR hold340/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06179_ _13851_/Q _13852_/Q _13853_/Q _13854_/Q VGND VGND VPWR VPWR _06179_/X sky130_fd_sc_hd__or4_1
Xhold351 hold351/A VGND VGND VPWR VPWR hold351/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold362 hold362/A VGND VGND VPWR VPWR hold362/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold373 hold373/A VGND VGND VPWR VPWR hold373/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold384 hold384/A VGND VGND VPWR VPWR hold384/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_131_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold395 hold395/A VGND VGND VPWR VPWR hold395/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09938_ _13493_/Q _13682_/Q _09946_/S VGND VGND VPWR VPWR _09939_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09869_ _13688_/Q _09865_/A _09868_/Y _09776_/X VGND VGND VPWR VPWR _13688_/D sky130_fd_sc_hd__o211a_1
XFILLER_100_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11900_ _11900_/A VGND VGND VPWR VPWR _14257_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12880_ _12881_/CLK _12880_/D hold1/X VGND VGND VPWR VPWR _12880_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _11831_/A VGND VGND VPWR VPWR _14107_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _14722_/CLK _14550_/D VGND VGND VPWR VPWR _14550_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11365_/X _14072_/Q _11766_/S VGND VGND VPWR VPWR _11763_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13698_/CLK hold287/X VGND VGND VPWR VPWR _13501_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10713_ _10713_/A VGND VGND VPWR VPWR _12934_/D sky130_fd_sc_hd__clkbuf_1
X_14481_ _14733_/CLK _14481_/D VGND VGND VPWR VPWR _14481_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _11693_/A VGND VGND VPWR VPWR _14028_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13432_ _14588_/CLK hold62/X VGND VGND VPWR VPWR _13432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10644_ _14411_/Q hold354/A VGND VGND VPWR VPWR _14362_/D sky130_fd_sc_hd__xor2_1
XFILLER_139_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10575_ _10575_/A _10575_/B VGND VGND VPWR VPWR _12671_/D sky130_fd_sc_hd__nand2_1
X_13363_ _13366_/CLK _13363_/D repeater56/X VGND VGND VPWR VPWR _13363_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12314_ _12314_/A VGND VGND VPWR VPWR _14572_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13294_ _13294_/CLK hold134/X VGND VGND VPWR VPWR _13294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12245_ _12245_/A VGND VGND VPWR VPWR _14538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12176_ _12176_/A VGND VGND VPWR VPWR _14499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11127_ _11127_/A _11084_/X VGND VGND VPWR VPWR _11127_/X sky130_fd_sc_hd__or2b_1
XFILLER_111_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11058_ _14604_/Q _14566_/Q _14497_/Q _14449_/Q _11044_/X _11045_/X VGND VGND VPWR
+ VPWR _11059_/A sky130_fd_sc_hd__mux4_1
XFILLER_49_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10009_ _10009_/A VGND VGND VPWR VPWR _12670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14748_ _14749_/CLK _14748_/D VGND VGND VPWR VPWR _14748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14679_ _14679_/CLK _14679_/D VGND VGND VPWR VPWR hold96/A sky130_fd_sc_hd__dfxtp_1
X_07220_ _14588_/Q _13116_/Q VGND VGND VPWR VPWR _07796_/A sky130_fd_sc_hd__xor2_1
XFILLER_149_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater60 hold2/X VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__buf_12
XFILLER_158_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07151_ _07151_/A _07151_/B VGND VGND VPWR VPWR _07152_/B sky130_fd_sc_hd__nand2_1
XFILLER_145_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06102_ _06102_/A VGND VGND VPWR VPWR _13941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07082_ _07082_/A _07082_/B VGND VGND VPWR VPWR _07126_/A sky130_fd_sc_hd__and2_1
XFILLER_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06033_ _06361_/A _12336_/C VGND VGND VPWR VPWR _14633_/D sky130_fd_sc_hd__nand2_1
XFILLER_113_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07984_ _06976_/X _07983_/X _07932_/X VGND VGND VPWR VPWR _13277_/D sky130_fd_sc_hd__a21o_1
XFILLER_101_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09723_ _09723_/A _09723_/B VGND VGND VPWR VPWR _09726_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06935_ _06935_/A _06934_/X VGND VGND VPWR VPWR _06951_/C sky130_fd_sc_hd__or2b_1
X_09654_ _09654_/A VGND VGND VPWR VPWR _12839_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06866_ _13013_/Q _07911_/B VGND VGND VPWR VPWR _06868_/A sky130_fd_sc_hd__nand2_1
XFILLER_103_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08605_ _08605_/A VGND VGND VPWR VPWR _08607_/B sky130_fd_sc_hd__inv_2
XFILLER_15_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06797_ _06793_/Y _06794_/X _06796_/X _06703_/X VGND VGND VPWR VPWR _13007_/D sky130_fd_sc_hd__a2bb2o_1
X_09585_ _13391_/Q _13589_/Q _09587_/S VGND VGND VPWR VPWR _09586_/A sky130_fd_sc_hd__mux2_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08536_ _08536_/A _08552_/B VGND VGND VPWR VPWR _09399_/B sky130_fd_sc_hd__xnor2_4
X_08467_ _14253_/Q _14251_/Q _08472_/A VGND VGND VPWR VPWR _08467_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07418_ _07428_/A _07298_/X _07329_/Y VGND VGND VPWR VPWR _07418_/X sky130_fd_sc_hd__o21ba_1
XFILLER_50_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08398_ _13095_/Q _13376_/Q _08406_/S VGND VGND VPWR VPWR _08399_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07349_ _07349_/A _07349_/B _07349_/C VGND VGND VPWR VPWR _07375_/B sky130_fd_sc_hd__and3_1
XFILLER_148_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10360_ _14211_/D VGND VGND VPWR VPWR _10432_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_109_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09019_ _09019_/A VGND VGND VPWR VPWR _12746_/D sky130_fd_sc_hd__clkbuf_1
X_10291_ _13522_/D VGND VGND VPWR VPWR _13469_/D sky130_fd_sc_hd__clkinv_2
X_12030_ _14682_/Q _12034_/B _12030_/C VGND VGND VPWR VPWR _12031_/A sky130_fd_sc_hd__and3_1
Xhold170 hold170/A VGND VGND VPWR VPWR hold170/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold181 hold181/A VGND VGND VPWR VPWR hold181/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold192 hold192/A VGND VGND VPWR VPWR hold192/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_160_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13981_ _14533_/CLK _13981_/D VGND VGND VPWR VPWR _13981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12932_ _13265_/CLK _12932_/D VGND VGND VPWR VPWR hold391/A sky130_fd_sc_hd__dfxtp_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _13700_/CLK _12863_/D VGND VGND VPWR VPWR hold127/A sky130_fd_sc_hd__dfxtp_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14602_/CLK _14602_/D VGND VGND VPWR VPWR _14602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11814_ _11814_/A VGND VGND VPWR VPWR _14099_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12794_ _14319_/CLK _12794_/D VGND VGND VPWR VPWR hold219/A sky130_fd_sc_hd__dfxtp_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _14533_/CLK _14533_/D VGND VGND VPWR VPWR _14533_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11323_/X _14064_/Q _11747_/S VGND VGND VPWR VPWR _11746_/A sky130_fd_sc_hd__mux2_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14464_ _14726_/CLK _14464_/D VGND VGND VPWR VPWR _14464_/Q sky130_fd_sc_hd__dfxtp_1
X_11676_ _14021_/Q _11475_/X _11678_/S VGND VGND VPWR VPWR _11677_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13415_ _14696_/CLK hold379/X VGND VGND VPWR VPWR _13415_/Q sky130_fd_sc_hd__dfxtp_1
X_10627_ _10627_/A _14394_/Q _14412_/Q VGND VGND VPWR VPWR _10627_/X sky130_fd_sc_hd__or3_1
XFILLER_155_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14395_ _14413_/CLK _14395_/D VGND VGND VPWR VPWR _14395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13346_ _14432_/CLK _13346_/D VGND VGND VPWR VPWR _13346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10558_ _10558_/A _10558_/B VGND VGND VPWR VPWR _10565_/A sky130_fd_sc_hd__or2_1
XFILLER_154_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13277_ _13283_/CLK _13277_/D repeater59/X VGND VGND VPWR VPWR _13277_/Q sky130_fd_sc_hd__dfrtp_2
X_10489_ _10490_/A _10490_/B _10490_/C VGND VGND VPWR VPWR _10498_/B sky130_fd_sc_hd__o21ai_1
X_12228_ _12278_/S VGND VGND VPWR VPWR _12237_/S sky130_fd_sc_hd__buf_2
XFILLER_97_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12159_ _14492_/Q _11962_/X _12161_/S VGND VGND VPWR VPWR _12160_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06720_ _06736_/A _06720_/B _06720_/C VGND VGND VPWR VPWR _06753_/A sky130_fd_sc_hd__and3_1
XFILLER_64_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06651_ _06841_/B _06645_/X _06646_/X _06648_/X _06674_/C _06745_/A VGND VGND VPWR
+ VPWR _06652_/D sky130_fd_sc_hd__mux4_2
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06582_ _06580_/X _06609_/B _06582_/C VGND VGND VPWR VPWR _06583_/A sky130_fd_sc_hd__and3b_1
X_09370_ _13589_/Q _09370_/B VGND VGND VPWR VPWR _09371_/B sky130_fd_sc_hd__nand2_1
XFILLER_91_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08321_ _13378_/Q _08325_/D _08298_/X VGND VGND VPWR VPWR _08322_/B sky130_fd_sc_hd__o21ai_1
X_08252_ _13366_/Q _08252_/B VGND VGND VPWR VPWR _08253_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07203_ _07163_/C _07203_/B _07203_/C VGND VGND VPWR VPWR _07207_/A sky130_fd_sc_hd__and3b_1
X_08183_ _08181_/X _08182_/Y _08180_/B _07326_/X VGND VGND VPWR VPWR _13359_/D sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_4_12_0_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR clkbuf_4_12_0_clk/X sky130_fd_sc_hd__clkbuf_2
X_07134_ _07133_/B _07134_/B VGND VGND VPWR VPWR _07135_/B sky130_fd_sc_hd__and2b_1
XFILLER_146_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07065_ _07119_/B _07086_/C _07141_/B hold425/A VGND VGND VPWR VPWR _07067_/A sky130_fd_sc_hd__a22oi_1
XFILLER_145_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06016_ hold173/A _13556_/Q _13557_/Q _06016_/D VGND VGND VPWR VPWR _06017_/D sky130_fd_sc_hd__or4_1
XFILLER_161_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07967_ _07970_/B _07966_/X _06930_/X VGND VGND VPWR VPWR _13274_/D sky130_fd_sc_hd__o21bai_1
XFILLER_102_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09706_ _13670_/Q _09707_/B VGND VGND VPWR VPWR _09725_/A sky130_fd_sc_hd__nor2_1
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06918_ _06919_/A _06919_/B _06924_/D VGND VGND VPWR VPWR _06918_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07898_ _07898_/A _07898_/B VGND VGND VPWR VPWR _07904_/B sky130_fd_sc_hd__and2_1
XFILLER_28_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09637_ _09637_/A VGND VGND VPWR VPWR _12831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06849_ _06871_/A _07895_/B _07895_/C VGND VGND VPWR VPWR _06849_/X sky130_fd_sc_hd__and3_1
XFILLER_130_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09568_ _13618_/Q _09569_/B VGND VGND VPWR VPWR _09568_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08519_ _08521_/A _08509_/B _08520_/C _08671_/A VGND VGND VPWR VPWR _08532_/B sky130_fd_sc_hd__a22o_1
XFILLER_70_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09499_ _09500_/A _09500_/B _09509_/C VGND VGND VPWR VPWR _09505_/B sky130_fd_sc_hd__a21o_1
XFILLER_23_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11530_ _11530_/A VGND VGND VPWR VPWR _13849_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11461_ _11461_/A VGND VGND VPWR VPWR _13822_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13200_ _13617_/CLK _13200_/D VGND VGND VPWR VPWR hold449/A sky130_fd_sc_hd__dfxtp_1
X_10412_ _10405_/A _10403_/X _10431_/A _10378_/A VGND VGND VPWR VPWR _10418_/B sky130_fd_sc_hd__o2bb2a_1
X_14180_ _14180_/CLK _14180_/D VGND VGND VPWR VPWR _14180_/Q sky130_fd_sc_hd__dfxtp_1
X_11392_ _13720_/Q _11394_/B VGND VGND VPWR VPWR _11393_/A sky130_fd_sc_hd__and2_1
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13131_ _13524_/CLK _13131_/D hold1/X VGND VGND VPWR VPWR _13131_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10343_ _14622_/Q _14623_/Q VGND VGND VPWR VPWR _10344_/B sky130_fd_sc_hd__and2_1
X_10274_ _12875_/Q _14326_/Q _14595_/Q VGND VGND VPWR VPWR _10275_/B sky130_fd_sc_hd__mux2_1
XFILLER_155_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13062_ _13587_/CLK _13062_/D VGND VGND VPWR VPWR hold298/A sky130_fd_sc_hd__dfxtp_1
XFILLER_140_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12013_ _12013_/A VGND VGND VPWR VPWR _12013_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13964_ _13964_/CLK _13964_/D VGND VGND VPWR VPWR _13964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12915_ _14697_/CLK _12915_/D VGND VGND VPWR VPWR hold238/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13895_ _14050_/CLK hold286/X VGND VGND VPWR VPWR _13895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ _13727_/CLK _12846_/D VGND VGND VPWR VPWR hold436/A sky130_fd_sc_hd__dfxtp_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _13565_/CLK _12777_/D VGND VGND VPWR VPWR hold151/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14608_/CLK _14516_/D VGND VGND VPWR VPWR _14516_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11728_ _11297_/X _14056_/Q _11736_/S VGND VGND VPWR VPWR _11729_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14447_ _14495_/CLK _14447_/D VGND VGND VPWR VPWR _14447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11659_ _14013_/Q _11446_/X _11667_/S VGND VGND VPWR VPWR _11660_/A sky130_fd_sc_hd__mux2_1
X_14378_ _14732_/CLK _14379_/Q VGND VGND VPWR VPWR hold520/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13329_ _14602_/CLK _13329_/D VGND VGND VPWR VPWR _13329_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_clk clkbuf_3_1_0_clk/A VGND VGND VPWR VPWR clkbuf_4_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_131_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08870_ _08870_/A _08870_/B VGND VGND VPWR VPWR _08914_/A sky130_fd_sc_hd__and2_1
XFILLER_85_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07821_ _13254_/Q _07821_/B VGND VGND VPWR VPWR _07821_/X sky130_fd_sc_hd__and2_1
XFILLER_84_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07752_ _07772_/D VGND VGND VPWR VPWR _07785_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06703_ _06859_/A VGND VGND VPWR VPWR _06703_/X sky130_fd_sc_hd__clkbuf_2
X_07683_ _07683_/A _07683_/B VGND VGND VPWR VPWR _07684_/B sky130_fd_sc_hd__xnor2_1
XFILLER_64_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09422_ _08577_/B _09421_/X _09422_/S VGND VGND VPWR VPWR _09423_/A sky130_fd_sc_hd__mux2_1
X_06634_ _13034_/Q _13039_/Q VGND VGND VPWR VPWR _06634_/X sky130_fd_sc_hd__and2b_1
X_09353_ _09353_/A VGND VGND VPWR VPWR _12802_/D sky130_fd_sc_hd__clkbuf_1
X_06565_ _12891_/Q _06565_/B VGND VGND VPWR VPWR _06566_/B sky130_fd_sc_hd__nor2_1
XFILLER_80_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08304_ _13372_/Q _08294_/A _08301_/D _13373_/Q VGND VGND VPWR VPWR _08305_/C sky130_fd_sc_hd__a31o_1
X_09284_ _13553_/Q _09284_/B VGND VGND VPWR VPWR _09285_/B sky130_fd_sc_hd__or2_1
X_06496_ _06496_/A VGND VGND VPWR VPWR _06500_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08235_ _08223_/Y _08214_/B _08222_/A _08211_/A VGND VGND VPWR VPWR _08236_/B sky130_fd_sc_hd__a211o_1
XFILLER_5_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08166_ _13358_/Q _08166_/B VGND VGND VPWR VPWR _08167_/B sky130_fd_sc_hd__or2_1
XFILLER_118_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07117_ _13115_/D VGND VGND VPWR VPWR _07190_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_08097_ _08097_/A VGND VGND VPWR VPWR _10781_/A sky130_fd_sc_hd__clkbuf_2
X_07048_ _07059_/B _07074_/B VGND VGND VPWR VPWR _07049_/B sky130_fd_sc_hd__nor2_1
XFILLER_133_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08999_ _08999_/A VGND VGND VPWR VPWR _14254_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10961_ _10932_/X _10957_/Y _10960_/Y _10946_/X VGND VGND VPWR VPWR _10962_/B sky130_fd_sc_hd__a211o_1
XFILLER_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12700_ _13314_/CLK _12700_/D VGND VGND VPWR VPWR hold74/A sky130_fd_sc_hd__dfxtp_1
X_13680_ _13680_/CLK _13680_/D repeater56/X VGND VGND VPWR VPWR _13680_/Q sky130_fd_sc_hd__dfrtp_1
X_10892_ _10892_/A VGND VGND VPWR VPWR _13204_/D sky130_fd_sc_hd__clkbuf_1
X_12631_ _14742_/Q _12631_/B _12631_/C VGND VGND VPWR VPWR _12635_/B sky130_fd_sc_hd__and3_1
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12562_ _11375_/X _14726_/Q _12562_/S VGND VGND VPWR VPWR _12563_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14301_ _14600_/CLK _14301_/D VGND VGND VPWR VPWR _14301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11513_ _12016_/A VGND VGND VPWR VPWR _11513_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12493_ _12493_/A VGND VGND VPWR VPWR _14676_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14232_ _14543_/CLK _14232_/D VGND VGND VPWR VPWR _14232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11444_ _13843_/D _11444_/B VGND VGND VPWR VPWR _11445_/A sky130_fd_sc_hd__and2_1
XFILLER_109_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14163_ _14209_/CLK _14163_/D VGND VGND VPWR VPWR hold419/A sky130_fd_sc_hd__dfxtp_1
X_11375_ _12025_/A VGND VGND VPWR VPWR _11375_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13114_ _14645_/CLK hold154/X VGND VGND VPWR VPWR _13114_/Q sky130_fd_sc_hd__dfxtp_1
X_10326_ _10330_/B _10326_/B VGND VGND VPWR VPWR _10327_/A sky130_fd_sc_hd__or2_1
XFILLER_3_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14094_ _14098_/CLK _14094_/D VGND VGND VPWR VPWR _14094_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _13528_/CLK _13045_/D VGND VGND VPWR VPWR hold305/A sky130_fd_sc_hd__dfxtp_1
X_10257_ _10252_/X _10256_/X _14555_/D VGND VGND VPWR VPWR _10258_/A sky130_fd_sc_hd__mux2_1
X_10188_ _10266_/S VGND VGND VPWR VPWR _14556_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_66_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13947_ _13964_/CLK _13947_/D VGND VGND VPWR VPWR _13947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13878_ _14657_/CLK hold232/X VGND VGND VPWR VPWR _13878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12829_ _13653_/CLK _12829_/D VGND VGND VPWR VPWR hold445/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06350_ _14406_/D _14407_/D _14408_/D _06350_/D VGND VGND VPWR VPWR _06351_/C sky130_fd_sc_hd__or4_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06281_ _13813_/Q _13797_/Q _06281_/S VGND VGND VPWR VPWR _06282_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_150_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _14713_/CLK sky130_fd_sc_hd__clkbuf_16
X_08020_ _13283_/Q _08020_/B VGND VGND VPWR VPWR _08020_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09971_ _09971_/A VGND VGND VPWR VPWR _12871_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08922_ _08921_/B _08922_/B VGND VGND VPWR VPWR _08923_/B sky130_fd_sc_hd__and2b_1
XFILLER_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08853_ _08907_/B _08874_/C _08929_/B _13516_/D VGND VGND VPWR VPWR _08855_/A sky130_fd_sc_hd__a22oi_1
XFILLER_69_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07804_ _13253_/Q _07804_/B _07804_/C VGND VGND VPWR VPWR _07806_/A sky130_fd_sc_hd__and3_1
XFILLER_85_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08784_ _09502_/A VGND VGND VPWR VPWR _08784_/X sky130_fd_sc_hd__buf_2
X_05996_ _06341_/S VGND VGND VPWR VPWR _06345_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_84_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07735_ _07735_/A _07735_/B _07735_/C VGND VGND VPWR VPWR _07737_/A sky130_fd_sc_hd__or3_1
XFILLER_26_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07666_ _13110_/Q _13111_/Q _13247_/D _14584_/Q VGND VGND VPWR VPWR _07696_/A sky130_fd_sc_hd__and4_1
X_09405_ _09405_/A VGND VGND VPWR VPWR _13595_/D sky130_fd_sc_hd__clkbuf_1
X_06617_ _12905_/Q _06616_/A _06609_/B VGND VGND VPWR VPWR _06617_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07597_ _13111_/Q VGND VGND VPWR VPWR _07645_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09336_ _09336_/A VGND VGND VPWR VPWR _12794_/D sky130_fd_sc_hd__clkbuf_1
X_06548_ _06548_/A VGND VGND VPWR VPWR _06548_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09267_ _09267_/A _09267_/B VGND VGND VPWR VPWR _09267_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_141_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _14208_/CLK sky130_fd_sc_hd__clkbuf_16
X_06479_ _06473_/B _06477_/Y _06530_/S VGND VGND VPWR VPWR _06480_/A sky130_fd_sc_hd__mux2_1
X_08218_ _09116_/S VGND VGND VPWR VPWR _08218_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_154_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09198_ _13539_/Q _07579_/B _09195_/Y VGND VGND VPWR VPWR _09205_/A sky130_fd_sc_hd__a21oi_1
XFILLER_153_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08149_ _13357_/Q _08150_/B VGND VGND VPWR VPWR _08169_/A sky130_fd_sc_hd__nor2_1
XFILLER_161_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11160_ _14611_/Q _14573_/Q _14504_/Q _14456_/Q _11115_/X _11116_/X VGND VGND VPWR
+ VPWR _11161_/A sky130_fd_sc_hd__mux4_1
XFILLER_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10111_ _14184_/Q _14176_/Q _10617_/A VGND VGND VPWR VPWR _10111_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11091_ _11162_/A VGND VGND VPWR VPWR _11091_/X sky130_fd_sc_hd__buf_2
XFILLER_0_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10042_ _13801_/Q _13785_/Q _13935_/D VGND VGND VPWR VPWR _10043_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__clkbuf_1
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold63 hold63/A VGND VGND VPWR VPWR hold63/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold74 hold74/A VGND VGND VPWR VPWR hold74/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold85 hold85/A VGND VGND VPWR VPWR hold85/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold96 hold96/A VGND VGND VPWR VPWR hold96/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_13801_ _13945_/CLK _13801_/D VGND VGND VPWR VPWR _13801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11993_ _11993_/A VGND VGND VPWR VPWR _14307_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13732_ _13805_/CLK hold341/X VGND VGND VPWR VPWR _13732_/Q sky130_fd_sc_hd__dfxtp_1
X_10944_ _10944_/A _10944_/B VGND VGND VPWR VPWR _10944_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13663_ _13666_/CLK _13663_/D VGND VGND VPWR VPWR _13663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10875_ _10875_/A VGND VGND VPWR VPWR _13196_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12614_ _12614_/A _12619_/B VGND VGND VPWR VPWR _12614_/Y sky130_fd_sc_hd__nor2_1
X_13594_ _13596_/CLK _13594_/D repeater56/X VGND VGND VPWR VPWR _13594_/Q sky130_fd_sc_hd__dfrtp_1
X_12545_ _12545_/A VGND VGND VPWR VPWR _12554_/S sky130_fd_sc_hd__buf_2
XFILLER_61_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_132_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _14196_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_157_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12476_ _14669_/Q _12019_/A _12480_/S VGND VGND VPWR VPWR _12477_/A sky130_fd_sc_hd__mux2_1
X_14215_ _14440_/CLK _14215_/D VGND VGND VPWR VPWR _14215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_5 _12261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11427_ _13736_/Q _11427_/B VGND VGND VPWR VPWR _11428_/A sky130_fd_sc_hd__and2_1
XFILLER_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14146_ _14294_/CLK hold400/X VGND VGND VPWR VPWR _14146_/Q sky130_fd_sc_hd__dfxtp_1
X_11358_ _13892_/Q _11362_/C _11357_/Y VGND VGND VPWR VPWR _12016_/A sky130_fd_sc_hd__a21oi_4
XFILLER_98_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10309_ _10310_/A _13513_/D VGND VGND VPWR VPWR _10309_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14077_ _14610_/CLK hold317/X VGND VGND VPWR VPWR hold229/A sky130_fd_sc_hd__dfxtp_1
XFILLER_112_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11289_ _13757_/Q _11288_/X _11295_/S VGND VGND VPWR VPWR _11290_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ _14275_/CLK _13028_/D repeater59/X VGND VGND VPWR VPWR _13028_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_67_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07520_ _13153_/Q _09206_/B VGND VGND VPWR VPWR _07530_/A sky130_fd_sc_hd__and2_1
XFILLER_19_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07451_ _13146_/Q _09188_/B VGND VGND VPWR VPWR _07452_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06402_ _10679_/A _06391_/A _06399_/X VGND VGND VPWR VPWR _06402_/Y sky130_fd_sc_hd__a21oi_1
X_07382_ _13139_/Q _07365_/X _07369_/X VGND VGND VPWR VPWR _07383_/B sky130_fd_sc_hd__a21bo_1
XFILLER_148_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09121_ _09114_/A _09134_/A _09119_/Y _09120_/Y VGND VGND VPWR VPWR _09122_/B sky130_fd_sc_hd__a31o_1
X_06333_ _14103_/Q _14087_/Q _06341_/S VGND VGND VPWR VPWR _06334_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_123_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _13698_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14756__67 VGND VGND VPWR VPWR _14756__67/HI data_o[30] sky130_fd_sc_hd__conb_1
X_06264_ _06262_/Y _06263_/X _13975_/D VGND VGND VPWR VPWR _06265_/A sky130_fd_sc_hd__mux2_1
X_09052_ _09052_/A VGND VGND VPWR VPWR _12761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08003_ _08003_/A _08003_/B VGND VGND VPWR VPWR _08013_/B sky130_fd_sc_hd__or2_1
XFILLER_135_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06195_ _14426_/Q VGND VGND VPWR VPWR _10194_/A sky130_fd_sc_hd__clkbuf_2
Xhold500 hold500/A VGND VGND VPWR VPWR hold500/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold511 hold511/A VGND VGND VPWR VPWR hold511/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09954_ _09954_/A VGND VGND VPWR VPWR _12863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08905_ _13432_/Q VGND VGND VPWR VPWR _08978_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _13694_/Q _09885_/B VGND VGND VPWR VPWR _09886_/A sky130_fd_sc_hd__and2_1
XFILLER_106_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08836_ _08847_/B _08862_/B VGND VGND VPWR VPWR _08837_/B sky130_fd_sc_hd__nor2_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08767_ _08767_/A _08767_/B VGND VGND VPWR VPWR _08768_/B sky130_fd_sc_hd__nand2_1
XFILLER_73_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05979_ _05979_/A _05979_/B VGND VGND VPWR VPWR _11576_/A sky130_fd_sc_hd__nand2_2
XFILLER_73_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07718_ _07738_/A _07718_/B VGND VGND VPWR VPWR _07718_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ _08698_/A _08693_/B VGND VGND VPWR VPWR _08704_/B sky130_fd_sc_hd__or2b_1
XFILLER_25_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07649_ _07649_/A _07649_/B VGND VGND VPWR VPWR _07651_/A sky130_fd_sc_hd__nor2_1
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10660_ _14337_/Q _14334_/Q _14338_/Q VGND VGND VPWR VPWR _10661_/C sky130_fd_sc_hd__a21o_1
XFILLER_41_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09319_ _13297_/Q _13535_/Q _09321_/S VGND VGND VPWR VPWR _09320_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_114_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _13617_/CLK sky130_fd_sc_hd__clkbuf_16
X_10591_ _13621_/Q _13472_/Q _13470_/Q _08464_/X VGND VGND VPWR VPWR _13621_/D sky130_fd_sc_hd__o31a_1
XFILLER_139_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12330_ _14580_/Q _12022_/X _12332_/S VGND VGND VPWR VPWR _12331_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12261_ _12261_/A VGND VGND VPWR VPWR _12270_/S sky130_fd_sc_hd__buf_2
X_14000_ _14724_/CLK _14000_/D VGND VGND VPWR VPWR _14000_/Q sky130_fd_sc_hd__dfxtp_1
X_11212_ _11212_/A _11155_/X VGND VGND VPWR VPWR _11212_/X sky130_fd_sc_hd__or2b_1
XFILLER_123_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12192_ _14507_/Q _12010_/X _12194_/S VGND VGND VPWR VPWR _12193_/A sky130_fd_sc_hd__mux2_1
Xoutput31 _13328_/Q VGND VGND VPWR VPWR data_o[10] sky130_fd_sc_hd__buf_2
XFILLER_1_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput42 _13338_/Q VGND VGND VPWR VPWR data_o[20] sky130_fd_sc_hd__buf_2
XFILLER_134_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput53 _13327_/Q VGND VGND VPWR VPWR data_o[9] sky130_fd_sc_hd__buf_2
X_11143_ _14610_/Q _14572_/Q _14503_/Q _14455_/Q _11115_/X _11116_/X VGND VGND VPWR
+ VPWR _11144_/A sky130_fd_sc_hd__mux4_1
XFILLER_122_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11074_ _14266_/Q _14657_/Q _13764_/Q _14712_/Q _11020_/X _11021_/X VGND VGND VPWR
+ VPWR _11075_/B sky130_fd_sc_hd__mux4_1
XFILLER_49_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10025_ _10034_/S VGND VGND VPWR VPWR _10032_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_63_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14764_ input28/X VGND VGND VPWR VPWR _14764_/X sky130_fd_sc_hd__clkbuf_1
X_11976_ _14302_/Q _11975_/X _11982_/S VGND VGND VPWR VPWR _11977_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13715_ _13799_/CLK hold43/X VGND VGND VPWR VPWR _13715_/Q sky130_fd_sc_hd__dfxtp_1
X_10927_ _14748_/Q VGND VGND VPWR VPWR _11166_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14695_ _14749_/CLK _14695_/D VGND VGND VPWR VPWR _14695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13646_ _14327_/CLK hold430/X VGND VGND VPWR VPWR _13646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10858_ _10858_/A VGND VGND VPWR VPWR _13188_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13577_ _14319_/CLK hold47/X VGND VGND VPWR VPWR _13577_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_105_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _13704_/CLK sky130_fd_sc_hd__clkbuf_16
X_10789_ _10789_/A VGND VGND VPWR VPWR _13057_/D sky130_fd_sc_hd__clkbuf_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12528_ _11304_/X _14710_/Q _12532_/S VGND VGND VPWR VPWR _12529_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12459_ _14661_/Q _14518_/Q _12461_/S VGND VGND VPWR VPWR _12460_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14129_ _14292_/CLK hold327/X VGND VGND VPWR VPWR hold301/A sky130_fd_sc_hd__dfxtp_1
XFILLER_113_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06951_ _06951_/A _06951_/B _06951_/C _06951_/D VGND VGND VPWR VPWR _06951_/Y sky130_fd_sc_hd__nor4_1
X_05902_ _13803_/Q _13804_/Q _13805_/Q _13806_/Q VGND VGND VPWR VPWR _05903_/C sky130_fd_sc_hd__or4_1
X_09670_ _13667_/Q _09883_/B VGND VGND VPWR VPWR _09671_/B sky130_fd_sc_hd__nand2_1
X_06882_ _06885_/A VGND VGND VPWR VPWR _07962_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_95_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08621_ _08621_/A _08621_/B _08621_/C VGND VGND VPWR VPWR _08630_/C sky130_fd_sc_hd__or3_1
XFILLER_54_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08552_ _08552_/A _08552_/B _08552_/C VGND VGND VPWR VPWR _08582_/B sky130_fd_sc_hd__and3_1
XFILLER_51_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07503_ _07503_/A _07503_/B VGND VGND VPWR VPWR _07532_/A sky130_fd_sc_hd__nand2_1
XFILLER_35_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08483_ _08682_/A VGND VGND VPWR VPWR _08733_/A sky130_fd_sc_hd__buf_2
X_07434_ _07434_/A _07438_/B VGND VGND VPWR VPWR _07434_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_149_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07365_ _09130_/B VGND VGND VPWR VPWR _07365_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09104_ _09098_/B _09103_/Y _09116_/S VGND VGND VPWR VPWR _09105_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06316_ _14189_/D _14190_/D _14191_/D _06316_/D VGND VGND VPWR VPWR _06316_/X sky130_fd_sc_hd__and4_1
X_07296_ _09098_/B _07294_/Y _09182_/A VGND VGND VPWR VPWR _07297_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09035_ _09035_/A VGND VGND VPWR VPWR _12753_/D sky130_fd_sc_hd__clkbuf_1
X_06247_ _14094_/Q _12678_/Q _06345_/S VGND VGND VPWR VPWR _06248_/A sky130_fd_sc_hd__mux2_1
Xhold330 hold330/A VGND VGND VPWR VPWR hold330/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06178_ _06178_/A VGND VGND VPWR VPWR _14176_/D sky130_fd_sc_hd__clkbuf_1
Xhold341 hold341/A VGND VGND VPWR VPWR hold341/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold352 hold352/A VGND VGND VPWR VPWR hold352/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold363 hold363/A VGND VGND VPWR VPWR hold363/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold374 hold374/A VGND VGND VPWR VPWR hold374/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold385 hold385/A VGND VGND VPWR VPWR hold385/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold396 hold396/A VGND VGND VPWR VPWR hold396/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_117_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09937_ _13700_/Q VGND VGND VPWR VPWR _09946_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_132_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _09868_/A VGND VGND VPWR VPWR _09868_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08819_ _08819_/A _08929_/A VGND VGND VPWR VPWR _08820_/B sky130_fd_sc_hd__nand2_1
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09799_ _09799_/A VGND VGND VPWR VPWR _13677_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _13585_/Q _11834_/B VGND VGND VPWR VPWR _11831_/A sky130_fd_sc_hd__and2_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11761_/A VGND VGND VPWR VPWR _14071_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13500_ _13700_/CLK hold277/X VGND VGND VPWR VPWR _13500_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _12891_/Q _10720_/B VGND VGND VPWR VPWR _10713_/A sky130_fd_sc_hd__and2_1
X_14480_ _14667_/CLK _14480_/D VGND VGND VPWR VPWR _14480_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _14028_/Q _11497_/X _11700_/S VGND VGND VPWR VPWR _11693_/A sky130_fd_sc_hd__mux2_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13431_ _14588_/CLK hold64/X VGND VGND VPWR VPWR _13431_/Q sky130_fd_sc_hd__dfxtp_1
X_10643_ _14165_/Q _10643_/B VGND VGND VPWR VPWR _14141_/D sky130_fd_sc_hd__xnor2_1
XFILLER_42_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13362_ _13362_/CLK _13362_/D repeater56/X VGND VGND VPWR VPWR _13362_/Q sky130_fd_sc_hd__dfrtp_1
X_10574_ _10574_/A VGND VGND VPWR VPWR _14439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12313_ _14572_/Q _11997_/X _12313_/S VGND VGND VPWR VPWR _12314_/A sky130_fd_sc_hd__mux2_1
X_13293_ _13294_/CLK hold248/X VGND VGND VPWR VPWR _13293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12244_ _11304_/X _14538_/Q _12248_/S VGND VGND VPWR VPWR _12245_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12175_ _14499_/Q _11984_/X _12183_/S VGND VGND VPWR VPWR _12176_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11126_ _14026_/Q _13992_/Q _13832_/Q _14544_/Q _11081_/X _11082_/X VGND VGND VPWR
+ VPWR _11127_/A sky130_fd_sc_hd__mux4_1
XFILLER_150_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11057_ _10991_/X _11054_/X _11056_/X _11015_/X VGND VGND VPWR VPWR _11057_/X sky130_fd_sc_hd__o211a_1
XFILLER_49_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10008_ _10007_/X _10004_/X _10008_/S VGND VGND VPWR VPWR _10009_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14747_ _14749_/CLK _14747_/D VGND VGND VPWR VPWR _14747_/Q sky130_fd_sc_hd__dfxtp_1
X_11959_ _14696_/Q VGND VGND VPWR VPWR _11959_/X sky130_fd_sc_hd__clkbuf_2
X_14678_ _14678_/CLK _14678_/D VGND VGND VPWR VPWR hold90/A sky130_fd_sc_hd__dfxtp_1
X_13629_ _14075_/CLK hold153/X VGND VGND VPWR VPWR _13629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07150_ _07150_/A _07150_/B VGND VGND VPWR VPWR _07152_/A sky130_fd_sc_hd__xnor2_2
XFILLER_146_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06101_ _13795_/Q _06105_/B VGND VGND VPWR VPWR _06102_/A sky130_fd_sc_hd__and2_1
XFILLER_157_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07081_ _07081_/A VGND VGND VPWR VPWR _13345_/D sky130_fd_sc_hd__clkbuf_1
X_06032_ _14642_/Q _14644_/Q _06032_/C VGND VGND VPWR VPWR _12336_/C sky130_fd_sc_hd__or3_1
XFILLER_145_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07983_ _07986_/B _07983_/B VGND VGND VPWR VPWR _07983_/X sky130_fd_sc_hd__xor2_1
XFILLER_86_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09722_ _13671_/Q _09722_/B VGND VGND VPWR VPWR _09723_/B sky130_fd_sc_hd__or2_1
X_06934_ _13019_/Q _06938_/B VGND VGND VPWR VPWR _06934_/X sky130_fd_sc_hd__or2_1
XFILLER_67_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09653_ _13422_/Q _13620_/Q _09653_/S VGND VGND VPWR VPWR _09654_/A sky130_fd_sc_hd__mux2_1
X_06865_ _07910_/B VGND VGND VPWR VPWR _07911_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08604_ _08464_/X _08601_/X _08603_/X VGND VGND VPWR VPWR _13445_/D sky130_fd_sc_hd__a21o_1
X_09584_ _09582_/Y _09583_/X _09493_/A VGND VGND VPWR VPWR _13620_/D sky130_fd_sc_hd__o21bai_1
X_06796_ _06796_/A _07863_/C VGND VGND VPWR VPWR _06796_/X sky130_fd_sc_hd__and2_1
XFILLER_36_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08535_ _08535_/A _08535_/B VGND VGND VPWR VPWR _08552_/B sky130_fd_sc_hd__and2_2
XFILLER_51_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08466_ _13473_/Q _14255_/Q _08472_/A VGND VGND VPWR VPWR _08645_/B sky130_fd_sc_hd__mux2_1
XFILLER_23_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07417_ _07338_/X _07367_/Y _07415_/C _07416_/X _07355_/A VGND VGND VPWR VPWR _07425_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_50_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08397_ _08397_/A VGND VGND VPWR VPWR _08406_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07348_ _07327_/X _07345_/X _07347_/X _07311_/A VGND VGND VPWR VPWR _07349_/C sky130_fd_sc_hd__o211a_1
XFILLER_6_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07279_ _07455_/A _09101_/B VGND VGND VPWR VPWR _07279_/X sky130_fd_sc_hd__and2_1
XFILLER_152_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09018_ _13210_/Q _13439_/Q _09018_/S VGND VGND VPWR VPWR _09019_/A sky130_fd_sc_hd__mux2_1
X_10290_ hold99/X VGND VGND VPWR VPWR _13165_/D sky130_fd_sc_hd__clkinv_2
XFILLER_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold160 hold160/A VGND VGND VPWR VPWR hold160/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold171 hold171/A VGND VGND VPWR VPWR hold171/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold182 hold182/A VGND VGND VPWR VPWR hold182/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_78_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold193 hold4/X VGND VGND VPWR VPWR hold193/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_160_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13980_ _14703_/CLK _13980_/D VGND VGND VPWR VPWR _13980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12931_ _13265_/CLK _12931_/D VGND VGND VPWR VPWR hold282/A sky130_fd_sc_hd__dfxtp_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ _13805_/CLK _12862_/D VGND VGND VPWR VPWR hold231/A sky130_fd_sc_hd__dfxtp_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _14712_/CLK _14601_/D VGND VGND VPWR VPWR _14601_/Q sky130_fd_sc_hd__dfxtp_1
X_11813_ _13577_/Q _11817_/B VGND VGND VPWR VPWR _11814_/A sky130_fd_sc_hd__and2_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _13574_/CLK _12793_/D VGND VGND VPWR VPWR hold269/A sky130_fd_sc_hd__dfxtp_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14725_/CLK _14532_/D VGND VGND VPWR VPWR _14532_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _11744_/A VGND VGND VPWR VPWR _14063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14463_ _14619_/CLK _14463_/D VGND VGND VPWR VPWR _14463_/Q sky130_fd_sc_hd__dfxtp_1
X_11675_ _11675_/A VGND VGND VPWR VPWR _14020_/D sky130_fd_sc_hd__clkbuf_1
X_13414_ _13617_/CLK hold362/X VGND VGND VPWR VPWR _13414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10626_ _10626_/A _10626_/B _10626_/C _10626_/D VGND VGND VPWR VPWR _10626_/X sky130_fd_sc_hd__or4_1
XFILLER_139_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14394_ _14413_/CLK _14394_/D VGND VGND VPWR VPWR _14394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13345_ _14432_/CLK _13345_/D VGND VGND VPWR VPWR _13345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10557_ _10557_/A _10557_/B _10557_/C VGND VGND VPWR VPWR _10558_/B sky130_fd_sc_hd__and3_1
XFILLER_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13276_ _13283_/CLK _13276_/D repeater59/X VGND VGND VPWR VPWR _13276_/Q sky130_fd_sc_hd__dfrtp_2
X_10488_ _10493_/A _10488_/B VGND VGND VPWR VPWR _10490_/C sky130_fd_sc_hd__xnor2_1
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12227_ _12261_/A VGND VGND VPWR VPWR _12278_/S sky130_fd_sc_hd__buf_2
XFILLER_142_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12158_ _12158_/A VGND VGND VPWR VPWR _14491_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11109_ _13329_/Q _11079_/X _11102_/X _11108_/Y VGND VGND VPWR VPWR _13329_/D sky130_fd_sc_hd__o22a_1
XFILLER_68_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12089_ _11365_/X _14462_/Q _12093_/S VGND VGND VPWR VPWR _12090_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06650_ _13039_/Q VGND VGND VPWR VPWR _06745_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06581_ _06574_/X _06584_/D _12894_/Q VGND VGND VPWR VPWR _06582_/C sky130_fd_sc_hd__a21o_1
XFILLER_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08320_ _13378_/Q _08325_/D VGND VGND VPWR VPWR _08322_/A sky130_fd_sc_hd__and2_1
X_08251_ _13366_/Q _08252_/B VGND VGND VPWR VPWR _08253_/A sky130_fd_sc_hd__and2_1
XFILLER_32_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07202_ _07178_/A _07205_/C _07197_/A VGND VGND VPWR VPWR _07208_/A sky130_fd_sc_hd__a21o_1
X_08182_ _08167_/A _08170_/X _08180_/Y VGND VGND VPWR VPWR _08182_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07133_ _07134_/B _07133_/B VGND VGND VPWR VPWR _07153_/B sky130_fd_sc_hd__and2b_1
XFILLER_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07064_ _07064_/A _07106_/A VGND VGND VPWR VPWR _07082_/A sky130_fd_sc_hd__nor2_1
XFILLER_145_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06015_ _13559_/Q _13560_/Q _13561_/Q _13562_/Q VGND VGND VPWR VPWR _06016_/D sky130_fd_sc_hd__or4_1
XFILLER_133_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07966_ _07957_/A _07961_/X _07972_/C _06836_/X VGND VGND VPWR VPWR _07966_/X sky130_fd_sc_hd__a31o_1
XFILLER_68_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09705_ _09702_/X _09704_/X _09758_/A VGND VGND VPWR VPWR _09707_/B sky130_fd_sc_hd__o21a_1
XFILLER_56_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06917_ _13017_/Q _06938_/B VGND VGND VPWR VPWR _06924_/D sky130_fd_sc_hd__xnor2_1
XFILLER_74_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07897_ _07905_/A _07904_/A VGND VGND VPWR VPWR _07917_/A sky130_fd_sc_hd__nor2_1
XFILLER_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_94_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _13722_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09636_ _13414_/Q _13612_/Q _09642_/S VGND VGND VPWR VPWR _09637_/A sky130_fd_sc_hd__mux2_1
X_06848_ _06851_/A _06857_/A _06851_/B VGND VGND VPWR VPWR _06848_/X sky130_fd_sc_hd__or3b_1
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09567_ _09565_/Y _09566_/X _09493_/A VGND VGND VPWR VPWR _13617_/D sky130_fd_sc_hd__o21bai_1
X_06779_ _06703_/X _06781_/B _06794_/B _06778_/Y VGND VGND VPWR VPWR _13006_/D sky130_fd_sc_hd__a22o_1
XFILLER_130_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08518_ _08427_/A _08635_/B _08444_/X _08445_/X _08473_/C _08544_/A VGND VGND VPWR
+ VPWR _08520_/C sky130_fd_sc_hd__mux4_1
X_09498_ _09505_/A _09498_/B VGND VGND VPWR VPWR _09509_/C sky130_fd_sc_hd__nand2_1
XFILLER_12_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08449_ _08635_/B _08444_/X _08445_/X _08446_/X _08473_/C _08544_/A VGND VGND VPWR
+ VPWR _08450_/D sky130_fd_sc_hd__mux4_2
XFILLER_12_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11460_ _13822_/Q _11459_/X _11463_/S VGND VGND VPWR VPWR _11461_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10411_ _10411_/A _10411_/B _10411_/C VGND VGND VPWR VPWR _10421_/B sky130_fd_sc_hd__and3_1
XFILLER_109_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11391_ _11391_/A VGND VGND VPWR VPWR _13788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13130_ _13294_/CLK hold500/X VGND VGND VPWR VPWR hold99/A sky130_fd_sc_hd__dfxtp_2
XFILLER_124_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10342_ _14622_/Q _14623_/Q VGND VGND VPWR VPWR _10348_/B sky130_fd_sc_hd__nor2_2
XFILLER_3_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13061_ _13587_/CLK _13061_/D VGND VGND VPWR VPWR hold297/A sky130_fd_sc_hd__dfxtp_1
X_10273_ _10593_/A _14323_/Q VGND VGND VPWR VPWR _12508_/B sky130_fd_sc_hd__and2b_1
XFILLER_3_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12012_ _12012_/A VGND VGND VPWR VPWR _14313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13963_ _13963_/CLK _13963_/D VGND VGND VPWR VPWR _13963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_85_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _13476_/CLK sky130_fd_sc_hd__clkbuf_16
X_12914_ _14696_/CLK _12914_/D VGND VGND VPWR VPWR hold311/A sky130_fd_sc_hd__dfxtp_1
X_13894_ _14209_/CLK hold225/X VGND VGND VPWR VPWR _13894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12845_ _13727_/CLK _12845_/D VGND VGND VPWR VPWR hold137/A sky130_fd_sc_hd__dfxtp_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _13565_/CLK _12776_/D VGND VGND VPWR VPWR hold174/A sky130_fd_sc_hd__dfxtp_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _11749_/A VGND VGND VPWR VPWR _11736_/S sky130_fd_sc_hd__clkbuf_2
X_14515_ _14608_/CLK _14515_/D VGND VGND VPWR VPWR _14515_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14446_ _14495_/CLK _14446_/D VGND VGND VPWR VPWR _14446_/Q sky130_fd_sc_hd__dfxtp_1
X_11658_ _11708_/S VGND VGND VPWR VPWR _11667_/S sky130_fd_sc_hd__buf_2
XFILLER_128_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10609_ _10032_/S _10606_/X _10607_/X _10608_/X _13934_/Q VGND VGND VPWR VPWR _13976_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14377_ _14536_/CLK hold520/X VGND VGND VPWR VPWR _14377_/Q sky130_fd_sc_hd__dfxtp_1
X_11589_ _13652_/Q _11591_/B VGND VGND VPWR VPWR _11590_/A sky130_fd_sc_hd__and2_1
X_13328_ _14602_/CLK _13328_/D VGND VGND VPWR VPWR _13328_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_127_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13259_ _13264_/CLK _13259_/D repeater59/X VGND VGND VPWR VPWR _13259_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07820_ _07833_/A _07820_/B VGND VGND VPWR VPWR _07823_/A sky130_fd_sc_hd__or2_1
XFILLER_57_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07751_ _07787_/A _07787_/B VGND VGND VPWR VPWR _07756_/A sky130_fd_sc_hd__xnor2_1
XFILLER_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_76_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _13362_/CLK sky130_fd_sc_hd__clkbuf_16
X_06702_ _06702_/A VGND VGND VPWR VPWR _13001_/D sky130_fd_sc_hd__clkbuf_1
X_07682_ _07713_/A _07713_/B VGND VGND VPWR VPWR _07683_/B sky130_fd_sc_hd__xnor2_1
XFILLER_53_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09421_ _09421_/A _09421_/B VGND VGND VPWR VPWR _09421_/X sky130_fd_sc_hd__xor2_1
XFILLER_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06633_ _13344_/Q _13342_/Q _06704_/S VGND VGND VPWR VPWR _06633_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09352_ _13312_/Q _13550_/Q _09354_/S VGND VGND VPWR VPWR _09353_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06564_ _12891_/Q _06565_/B VGND VGND VPWR VPWR _06566_/A sky130_fd_sc_hd__and2_1
XFILLER_21_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08303_ _08303_/A VGND VGND VPWR VPWR _09084_/A sky130_fd_sc_hd__buf_4
X_09283_ _13553_/Q _09284_/B VGND VGND VPWR VPWR _09285_/A sky130_fd_sc_hd__nand2_1
XFILLER_100_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06495_ _06502_/A _10349_/A _06495_/C VGND VGND VPWR VPWR _06496_/A sky130_fd_sc_hd__and3_1
XFILLER_139_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08234_ _08234_/A VGND VGND VPWR VPWR _08236_/A sky130_fd_sc_hd__inv_2
XFILLER_147_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08165_ _13358_/Q _08166_/B VGND VGND VPWR VPWR _08167_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07116_ hold154/A VGND VGND VPWR VPWR _07190_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08096_ _08096_/A VGND VGND VPWR VPWR _12707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07047_ _07044_/Y _07074_/A _14634_/Q _07163_/A VGND VGND VPWR VPWR _07074_/B sky130_fd_sc_hd__and4bb_1
XFILLER_0_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08998_ _08986_/Y _08997_/Y _09006_/S VGND VGND VPWR VPWR _08999_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07949_ _07949_/A _07949_/B _07949_/C _07949_/D VGND VGND VPWR VPWR _07973_/A sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_67_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _13532_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_141_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10960_ _10960_/A _10960_/B VGND VGND VPWR VPWR _10960_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09619_ _09619_/A VGND VGND VPWR VPWR _12823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10891_ _13162_/Q _10891_/B VGND VGND VPWR VPWR _10892_/A sky130_fd_sc_hd__and2_1
XFILLER_34_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12630_ _12631_/B _12631_/C _12629_/Y VGND VGND VPWR VPWR _14741_/D sky130_fd_sc_hd__a21oi_1
XFILLER_71_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12561_ _12561_/A VGND VGND VPWR VPWR _14725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14300_ _14495_/CLK _14300_/D VGND VGND VPWR VPWR _14300_/Q sky130_fd_sc_hd__dfxtp_1
X_11512_ _11512_/A VGND VGND VPWR VPWR _13838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12492_ _12496_/A _12496_/B input13/X VGND VGND VPWR VPWR _12493_/A sky130_fd_sc_hd__and3_1
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14231_ _14543_/CLK _14231_/D VGND VGND VPWR VPWR _14231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11443_ _11443_/A VGND VGND VPWR VPWR _13812_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14162_ _14209_/CLK hold199/X VGND VGND VPWR VPWR _14162_/Q sky130_fd_sc_hd__dfxtp_1
X_11374_ _11373_/Y _13925_/Q _13878_/Q VGND VGND VPWR VPWR _12025_/A sky130_fd_sc_hd__a21o_4
XFILLER_109_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13113_ _14645_/CLK hold177/X VGND VGND VPWR VPWR _13113_/Q sky130_fd_sc_hd__dfxtp_1
X_10325_ _13747_/Q _13748_/Q VGND VGND VPWR VPWR _10326_/B sky130_fd_sc_hd__and2_1
X_14093_ _14319_/CLK _14093_/D VGND VGND VPWR VPWR _14093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _13528_/CLK _13044_/D VGND VGND VPWR VPWR hold294/A sky130_fd_sc_hd__dfxtp_1
X_10256_ _10247_/X _10255_/X _14556_/D VGND VGND VPWR VPWR _10256_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10187_ _10226_/A _14360_/Q VGND VGND VPWR VPWR _10266_/S sky130_fd_sc_hd__xor2_2
XFILLER_66_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_58_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _13666_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_11_0_clk clkbuf_3_5_0_clk/X VGND VGND VPWR VPWR clkbuf_4_11_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13946_ _13964_/CLK _13946_/D VGND VGND VPWR VPWR _13946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13877_ _14656_/CLK _13877_/D VGND VGND VPWR VPWR _13877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12828_ _13653_/CLK _12828_/D VGND VGND VPWR VPWR hold325/A sky130_fd_sc_hd__dfxtp_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _13602_/CLK _12759_/D VGND VGND VPWR VPWR hold110/A sky130_fd_sc_hd__dfxtp_1
XFILLER_148_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06280_ _06280_/A VGND VGND VPWR VPWR _13958_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14429_ _14643_/CLK _14429_/D VGND VGND VPWR VPWR _14429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09970_ _13508_/Q _13697_/Q _09974_/S VGND VGND VPWR VPWR _09971_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08921_ _08922_/B _08921_/B VGND VGND VPWR VPWR _08941_/B sky130_fd_sc_hd__and2b_1
XFILLER_115_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08852_ _08852_/A _08894_/A VGND VGND VPWR VPWR _08870_/A sky130_fd_sc_hd__nor2_1
XFILLER_29_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07803_ _07807_/B _07803_/B VGND VGND VPWR VPWR _13252_/D sky130_fd_sc_hd__xnor2_1
XFILLER_85_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08783_ _08706_/X _08781_/Y _08782_/X _08764_/X VGND VGND VPWR VPWR _13464_/D sky130_fd_sc_hd__a31o_1
XFILLER_84_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05995_ _06231_/A VGND VGND VPWR VPWR _06341_/S sky130_fd_sc_hd__inv_2
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_49_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _13351_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07734_ _07734_/A _07734_/B VGND VGND VPWR VPWR _07735_/C sky130_fd_sc_hd__xnor2_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07665_ _13111_/Q _13247_/D _14584_/Q _07645_/A VGND VGND VPWR VPWR _07665_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_53_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09404_ _09417_/B _09403_/X _09404_/S VGND VGND VPWR VPWR _09405_/A sky130_fd_sc_hd__mux2_1
X_06616_ _06616_/A _06616_/B VGND VGND VPWR VPWR _12904_/D sky130_fd_sc_hd__nor2_1
XFILLER_111_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07596_ _13244_/D VGND VGND VPWR VPWR _07701_/A sky130_fd_sc_hd__clkbuf_2
X_09335_ _13304_/Q _13542_/Q _09343_/S VGND VGND VPWR VPWR _09336_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06547_ _06547_/A _06547_/B VGND VGND VPWR VPWR _06550_/A sky130_fd_sc_hd__nor2_1
XFILLER_139_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09266_ _07239_/X _09265_/Y _07486_/X VGND VGND VPWR VPWR _13550_/D sky130_fd_sc_hd__a21o_1
X_06478_ _12910_/Q VGND VGND VPWR VPWR _06530_/S sky130_fd_sc_hd__buf_2
X_08217_ _13165_/Q VGND VGND VPWR VPWR _09116_/S sky130_fd_sc_hd__buf_2
X_09197_ _09195_/Y _09196_/X _07526_/X VGND VGND VPWR VPWR _13539_/D sky130_fd_sc_hd__o21bai_1
XFILLER_147_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08148_ _08145_/X _08147_/X _08199_/A VGND VGND VPWR VPWR _08150_/B sky130_fd_sc_hd__o21a_1
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08079_ _08079_/A VGND VGND VPWR VPWR _12699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10110_ _10110_/A VGND VGND VPWR VPWR _10617_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11090_ _11090_/A VGND VGND VPWR VPWR _11090_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10041_ _10041_/A VGND VGND VPWR VPWR _13946_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__buf_4
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold64 hold64/A VGND VGND VPWR VPWR hold64/X sky130_fd_sc_hd__clkbuf_2
Xhold75 hold75/A VGND VGND VPWR VPWR hold75/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold86 hold86/A VGND VGND VPWR VPWR hold86/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_13800_ _13945_/CLK _13800_/D VGND VGND VPWR VPWR _13800_/Q sky130_fd_sc_hd__dfxtp_1
Xhold97 hold97/A VGND VGND VPWR VPWR hold97/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_11992_ _14307_/Q _11991_/X _11998_/S VGND VGND VPWR VPWR _11993_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10943_ _14257_/Q _14648_/Q _13755_/Q _14703_/Q _10940_/X _10942_/X VGND VGND VPWR
+ VPWR _10944_/B sky130_fd_sc_hd__mux4_1
X_13731_ _13805_/CLK hold319/X VGND VGND VPWR VPWR _13731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_0_0_clk clkbuf_3_1_0_clk/A VGND VGND VPWR VPWR clkbuf_4_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_10874_ _13154_/Q _10874_/B VGND VGND VPWR VPWR _10875_/A sky130_fd_sc_hd__and2_1
X_13662_ _13666_/CLK _13662_/D VGND VGND VPWR VPWR _13662_/Q sky130_fd_sc_hd__dfxtp_1
X_12613_ _14734_/Q _12611_/A _12612_/Y VGND VGND VPWR VPWR _14734_/D sky130_fd_sc_hd__o21a_1
X_13593_ _13593_/CLK _13593_/D repeater56/X VGND VGND VPWR VPWR _13593_/Q sky130_fd_sc_hd__dfrtp_1
X_12544_ _12544_/A VGND VGND VPWR VPWR _14717_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12475_ _12475_/A VGND VGND VPWR VPWR _14668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14214_ _14440_/CLK _14214_/D VGND VGND VPWR VPWR _14214_/Q sky130_fd_sc_hd__dfxtp_1
X_11426_ _11426_/A VGND VGND VPWR VPWR _13804_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_6 _12261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14145_ _14159_/CLK _14145_/D VGND VGND VPWR VPWR _14145_/Q sky130_fd_sc_hd__dfxtp_1
X_11357_ _13892_/Q _11362_/C _11353_/B VGND VGND VPWR VPWR _11357_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_153_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10308_ _10304_/A _13512_/D _10307_/A VGND VGND VPWR VPWR _10312_/A sky130_fd_sc_hd__a21oi_1
X_14076_ _14610_/CLK hold229/X VGND VGND VPWR VPWR _14076_/Q sky130_fd_sc_hd__dfxtp_1
X_11288_ _14696_/Q VGND VGND VPWR VPWR _11288_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_141_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ _13027_/CLK _13027_/D repeater59/X VGND VGND VPWR VPWR _13027_/Q sky130_fd_sc_hd__dfrtp_1
X_10239_ _14526_/D _10238_/X _10266_/S VGND VGND VPWR VPWR _10240_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13929_ _14179_/CLK hold498/X VGND VGND VPWR VPWR _13929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07450_ _07450_/A VGND VGND VPWR VPWR _09188_/B sky130_fd_sc_hd__clkbuf_2
X_06401_ _10679_/A _06391_/A _06399_/X _06500_/A VGND VGND VPWR VPWR _06401_/X sky130_fd_sc_hd__a31o_1
X_07381_ _07381_/A _07415_/A VGND VGND VPWR VPWR _07416_/B sky130_fd_sc_hd__or2_1
X_09120_ _13528_/Q _09120_/B VGND VGND VPWR VPWR _09120_/Y sky130_fd_sc_hd__nor2_1
X_06332_ _06332_/A VGND VGND VPWR VPWR _14401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09051_ _13225_/Q _13454_/Q _09051_/S VGND VGND VPWR VPWR _09052_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06263_ hold498/A _13974_/D VGND VGND VPWR VPWR _06263_/X sky130_fd_sc_hd__and2_1
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08002_ _13280_/Q _08002_/B VGND VGND VPWR VPWR _08003_/B sky130_fd_sc_hd__nor2_1
XFILLER_163_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06194_ _06194_/A VGND VGND VPWR VPWR _14366_/D sky130_fd_sc_hd__clkbuf_1
Xhold501 hold501/A VGND VGND VPWR VPWR hold501/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold512 hold512/A VGND VGND VPWR VPWR hold512/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09953_ _13500_/Q _13689_/Q _09957_/S VGND VGND VPWR VPWR _09954_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08904_ _13431_/Q VGND VGND VPWR VPWR _08978_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _09884_/A VGND VGND VPWR VPWR _13693_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08835_ _08832_/Y _08862_/A _13515_/D _08951_/A VGND VGND VPWR VPWR _08862_/B sky130_fd_sc_hd__and4bb_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08766_ _13462_/Q _09555_/B VGND VGND VPWR VPWR _08770_/B sky130_fd_sc_hd__xnor2_1
X_05978_ _05965_/X _05966_/X _05970_/X _05977_/Y VGND VGND VPWR VPWR _05979_/B sky130_fd_sc_hd__a31o_1
XFILLER_122_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07717_ _07735_/B _07717_/B VGND VGND VPWR VPWR _07718_/B sky130_fd_sc_hd__or2_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08697_ _08617_/X _08694_/X _08695_/Y _08696_/X VGND VGND VPWR VPWR _13452_/D sky130_fd_sc_hd__a31o_1
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07648_ _13244_/D _13245_/D _07668_/C _13113_/Q VGND VGND VPWR VPWR _07649_/B sky130_fd_sc_hd__and4_1
XFILLER_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07579_ _13161_/Q _07579_/B VGND VGND VPWR VPWR _07581_/A sky130_fd_sc_hd__and2_1
XFILLER_22_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09318_ _09318_/A VGND VGND VPWR VPWR _12786_/D sky130_fd_sc_hd__clkbuf_1
X_10590_ _13555_/Q _13168_/Q hold487/A _07343_/X VGND VGND VPWR VPWR _13555_/D sky130_fd_sc_hd__o31a_1
X_09249_ _08218_/X _09247_/Y _09248_/X _09215_/X VGND VGND VPWR VPWR _13547_/D sky130_fd_sc_hd__a31o_1
XFILLER_154_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12260_ _12260_/A VGND VGND VPWR VPWR _14545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11211_ _14032_/Q _13998_/Q _13838_/Q _14550_/Q _11152_/X _11153_/X VGND VGND VPWR
+ VPWR _11212_/A sky130_fd_sc_hd__mux4_1
XFILLER_147_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12191_ _12191_/A VGND VGND VPWR VPWR _14506_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput32 _13329_/Q VGND VGND VPWR VPWR data_o[11] sky130_fd_sc_hd__buf_2
XFILLER_135_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput43 _13339_/Q VGND VGND VPWR VPWR data_o[21] sky130_fd_sc_hd__buf_2
X_11142_ _11136_/X _11139_/X _11141_/X _11086_/X VGND VGND VPWR VPWR _11142_/X sky130_fd_sc_hd__o211a_1
XFILLER_150_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput54 _14764_/X VGND VGND VPWR VPWR rtr_o sky130_fd_sc_hd__buf_2
XFILLER_150_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11073_ _11073_/A VGND VGND VPWR VPWR _11073_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10024_ _13952_/Q _13944_/Q _10607_/A VGND VGND VPWR VPWR _10024_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11975_ _14701_/Q VGND VGND VPWR VPWR _11975_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13714_ _13727_/CLK hold414/X VGND VGND VPWR VPWR _13714_/Q sky130_fd_sc_hd__dfxtp_1
X_10926_ _10926_/A _10925_/X VGND VGND VPWR VPWR _10926_/X sky130_fd_sc_hd__or2b_1
X_14694_ _14737_/CLK hold513/X VGND VGND VPWR VPWR _14694_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13645_ _14327_/CLK hold135/X VGND VGND VPWR VPWR _13645_/Q sky130_fd_sc_hd__dfxtp_1
X_10857_ _13146_/Q _10863_/B VGND VGND VPWR VPWR _10858_/A sky130_fd_sc_hd__and2_1
XFILLER_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13576_ _14319_/CLK hold55/X VGND VGND VPWR VPWR _13576_/Q sky130_fd_sc_hd__dfxtp_1
X_10788_ _13015_/Q _10790_/B VGND VGND VPWR VPWR _10789_/A sky130_fd_sc_hd__and2_1
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12527_ _12527_/A VGND VGND VPWR VPWR _14709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12458_ _12458_/A VGND VGND VPWR VPWR _14660_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11409_ _11409_/A VGND VGND VPWR VPWR _13796_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12389_ _12389_/A VGND VGND VPWR VPWR _14616_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14128_ _14159_/CLK hold395/X VGND VGND VPWR VPWR hold308/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06950_ _06950_/A _06950_/B VGND VGND VPWR VPWR _06951_/D sky130_fd_sc_hd__nand2_1
X_14059_ _14539_/CLK _14059_/D VGND VGND VPWR VPWR _14059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05901_ _13807_/Q _13808_/Q _13809_/Q _13810_/Q VGND VGND VPWR VPWR _05903_/B sky130_fd_sc_hd__or4_1
X_06881_ _06881_/A _06881_/B _06881_/C VGND VGND VPWR VPWR _06885_/A sky130_fd_sc_hd__and3_1
XFILLER_95_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08620_ _08620_/A _08620_/B _08620_/C VGND VGND VPWR VPWR _08621_/C sky130_fd_sc_hd__or3_1
XFILLER_39_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08551_ _08544_/X _08657_/B _08550_/X _08535_/A VGND VGND VPWR VPWR _08552_/C sky130_fd_sc_hd__o211a_1
XFILLER_82_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07502_ _13151_/Q _09212_/B VGND VGND VPWR VPWR _07503_/B sky130_fd_sc_hd__or2_1
X_08482_ _13469_/Q VGND VGND VPWR VPWR _08682_/A sky130_fd_sc_hd__inv_2
X_07433_ _13143_/Q _09163_/B _07424_/X VGND VGND VPWR VPWR _07438_/B sky130_fd_sc_hd__a21bo_1
XFILLER_149_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07364_ _07364_/A _07364_/B VGND VGND VPWR VPWR _09130_/B sky130_fd_sc_hd__xnor2_4
X_09103_ _09103_/A _09103_/B VGND VGND VPWR VPWR _09103_/Y sky130_fd_sc_hd__xnor2_1
X_06315_ hold199/A _14184_/D _14185_/D _14188_/D VGND VGND VPWR VPWR _06316_/D sky130_fd_sc_hd__and4_1
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07295_ _13165_/Q VGND VGND VPWR VPWR _09182_/A sky130_fd_sc_hd__buf_2
XFILLER_148_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09034_ _13217_/Q _13446_/Q _09040_/S VGND VGND VPWR VPWR _09035_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06246_ _06246_/A VGND VGND VPWR VPWR _14392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold320 hold320/A VGND VGND VPWR VPWR hold320/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold331 hold331/A VGND VGND VPWR VPWR hold331/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06177_ _13862_/Q _12679_/Q _06313_/S VGND VGND VPWR VPWR _06178_/A sky130_fd_sc_hd__mux2_1
Xhold342 hold342/A VGND VGND VPWR VPWR hold342/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold353 hold353/A VGND VGND VPWR VPWR hold353/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold364 hold364/A VGND VGND VPWR VPWR hold364/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold375 hold375/A VGND VGND VPWR VPWR hold375/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold386 hold386/A VGND VGND VPWR VPWR hold386/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold397 hold397/A VGND VGND VPWR VPWR hold397/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_120_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09936_ _09936_/A VGND VGND VPWR VPWR _12855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _09870_/B _09873_/D VGND VGND VPWR VPWR _09868_/A sky130_fd_sc_hd__and2_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08818_ _08874_/C VGND VGND VPWR VPWR _08929_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09798_ _09791_/B _09796_/Y _09834_/S VGND VGND VPWR VPWR _09799_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08749_ _08758_/A _08757_/A _08633_/A VGND VGND VPWR VPWR _08749_/X sky130_fd_sc_hd__o21a_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _11359_/X _14071_/Q _11766_/S VGND VGND VPWR VPWR _11761_/A sky130_fd_sc_hd__mux2_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _13031_/D VGND VGND VPWR VPWR _10720_/B sky130_fd_sc_hd__clkbuf_1
X_11691_ _11691_/A VGND VGND VPWR VPWR _11700_/S sky130_fd_sc_hd__buf_2
XFILLER_41_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13430_ _14588_/CLK hold79/X VGND VGND VPWR VPWR _13430_/Q sky130_fd_sc_hd__dfxtp_1
X_10642_ _14194_/Q _14197_/Q _14168_/Q VGND VGND VPWR VPWR _10643_/B sky130_fd_sc_hd__o21ai_1
XFILLER_41_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13361_ _13434_/CLK _13361_/D repeater56/X VGND VGND VPWR VPWR _13361_/Q sky130_fd_sc_hd__dfrtp_1
X_10573_ _10557_/C _10575_/B _10573_/C VGND VGND VPWR VPWR _10574_/A sky130_fd_sc_hd__and3b_1
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12312_ _12312_/A VGND VGND VPWR VPWR _14571_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13292_ _13296_/CLK hold307/X VGND VGND VPWR VPWR _13292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12243_ _12243_/A VGND VGND VPWR VPWR _14537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12174_ _12185_/A VGND VGND VPWR VPWR _12183_/S sky130_fd_sc_hd__buf_2
X_11125_ _14308_/Q _14478_/Q _14234_/Q _14064_/Q _11066_/X _11067_/X VGND VGND VPWR
+ VPWR _11125_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11056_ _11056_/A _11013_/X VGND VGND VPWR VPWR _11056_/X sky130_fd_sc_hd__or2b_1
XFILLER_67_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10007_ _13388_/Q _14627_/Q _10636_/A VGND VGND VPWR VPWR _10007_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14746_ _14746_/CLK _14746_/D VGND VGND VPWR VPWR _14746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11958_ _11958_/A VGND VGND VPWR VPWR _14296_/D sky130_fd_sc_hd__clkbuf_1
X_10909_ _12590_/A VGND VGND VPWR VPWR _11262_/A sky130_fd_sc_hd__buf_2
X_14677_ _14688_/CLK _14677_/D VGND VGND VPWR VPWR hold336/A sky130_fd_sc_hd__dfxtp_1
X_11889_ _11889_/A VGND VGND VPWR VPWR _14241_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13628_ _13635_/CLK hold406/X VGND VGND VPWR VPWR _13628_/Q sky130_fd_sc_hd__dfxtp_1
X_13559_ _13565_/CLK hold462/X VGND VGND VPWR VPWR _13559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06100_ _06100_/A VGND VGND VPWR VPWR _13940_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07080_ _07055_/Y _07079_/Y _10647_/A VGND VGND VPWR VPWR _07081_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06031_ _14645_/Q _14641_/Q _14643_/Q VGND VGND VPWR VPWR _06032_/C sky130_fd_sc_hd__or3_1
XFILLER_161_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07982_ _13276_/Q _08020_/B _07987_/A _07986_/A VGND VGND VPWR VPWR _07983_/B sky130_fd_sc_hd__a22o_1
X_06933_ _13019_/Q _06938_/B VGND VGND VPWR VPWR _06935_/A sky130_fd_sc_hd__and2_1
X_09721_ _13671_/Q _09722_/B VGND VGND VPWR VPWR _09723_/A sky130_fd_sc_hd__nand2_1
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09652_ _09652_/A VGND VGND VPWR VPWR _12838_/D sky130_fd_sc_hd__clkbuf_1
X_06864_ _06796_/A _06800_/B _06813_/C _06863_/X _06769_/B VGND VGND VPWR VPWR _07910_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_94_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08603_ _08642_/A _09438_/B VGND VGND VPWR VPWR _08603_/X sky130_fd_sc_hd__and2_1
X_09583_ _09577_/A _09578_/X _09581_/Y _08642_/A VGND VGND VPWR VPWR _09583_/X sky130_fd_sc_hd__a31o_1
XFILLER_82_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06795_ _07863_/B VGND VGND VPWR VPWR _06796_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08534_ _08427_/A _08645_/B _08467_/X _08471_/X _08579_/S _08544_/A VGND VGND VPWR
+ VPWR _08535_/B sky130_fd_sc_hd__mux4_1
XFILLER_36_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08465_ _08457_/B _08459_/B _08457_/A VGND VGND VPWR VPWR _08481_/A sky130_fd_sc_hd__o21ba_1
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07416_ _07416_/A _07416_/B VGND VGND VPWR VPWR _07416_/X sky130_fd_sc_hd__or2_1
X_08396_ _08396_/A VGND VGND VPWR VPWR _12730_/D sky130_fd_sc_hd__clkbuf_1
X_07347_ _07387_/A _07347_/B VGND VGND VPWR VPWR _07347_/X sky130_fd_sc_hd__or2_1
XFILLER_137_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07278_ _08157_/A VGND VGND VPWR VPWR _07455_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_164_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09017_ _09017_/A VGND VGND VPWR VPWR _12745_/D sky130_fd_sc_hd__clkbuf_1
X_06229_ _14415_/D _14416_/D VGND VGND VPWR VPWR _06230_/A sky130_fd_sc_hd__or2_1
XFILLER_152_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold150 input14/X VGND VGND VPWR VPWR hold150/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold161 hold161/A VGND VGND VPWR VPWR hold161/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold172 hold172/A VGND VGND VPWR VPWR hold172/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_160_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold183 hold183/A VGND VGND VPWR VPWR hold183/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold194 hold194/A VGND VGND VPWR VPWR hold194/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09919_ _09919_/A VGND VGND VPWR VPWR _12847_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12930_ _12930_/CLK _12930_/D VGND VGND VPWR VPWR hold112/A sky130_fd_sc_hd__dfxtp_1
XFILLER_59_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _13805_/CLK _12861_/D VGND VGND VPWR VPWR hold291/A sky130_fd_sc_hd__dfxtp_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _14600_/CLK _14600_/D VGND VGND VPWR VPWR _14600_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _11812_/A VGND VGND VPWR VPWR _14098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _13574_/CLK _12792_/D VGND VGND VPWR VPWR hold167/A sky130_fd_sc_hd__dfxtp_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _14533_/CLK _14531_/D VGND VGND VPWR VPWR _14531_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11320_/X _14063_/Q _11747_/S VGND VGND VPWR VPWR _11744_/A sky130_fd_sc_hd__mux2_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14462_ _14726_/CLK _14462_/D VGND VGND VPWR VPWR _14462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _14020_/Q _11472_/X _11678_/S VGND VGND VPWR VPWR _11675_/A sky130_fd_sc_hd__mux2_1
X_13413_ _13617_/CLK hold492/X VGND VGND VPWR VPWR _13413_/Q sky130_fd_sc_hd__dfxtp_1
X_10625_ _10623_/X _10624_/X hold28/X VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__o21a_1
X_14393_ _14410_/CLK _14393_/D VGND VGND VPWR VPWR _14393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13344_ _14432_/CLK _13344_/D VGND VGND VPWR VPWR _13344_/Q sky130_fd_sc_hd__dfxtp_1
X_10556_ _10557_/A _10573_/C _10557_/C VGND VGND VPWR VPWR _10558_/A sky130_fd_sc_hd__a21oi_1
XFILLER_127_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10487_ _10444_/B _10501_/C _10456_/C _10476_/A _10474_/A VGND VGND VPWR VPWR _10488_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_6_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13275_ _13283_/CLK _13275_/D repeater59/X VGND VGND VPWR VPWR _13275_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12226_ _12226_/A _12041_/C VGND VGND VPWR VPWR _12261_/A sky130_fd_sc_hd__or2b_4
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12157_ _14491_/Q _11959_/X _12161_/S VGND VGND VPWR VPWR _12158_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11108_ _11108_/A _11108_/B VGND VGND VPWR VPWR _11108_/Y sky130_fd_sc_hd__nand2_1
X_12088_ _12088_/A VGND VGND VPWR VPWR _14461_/D sky130_fd_sc_hd__clkbuf_1
X_11039_ _14302_/Q _14472_/Q _14228_/Q _14058_/Q _10993_/X _10995_/X VGND VGND VPWR
+ VPWR _11039_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06580_ _12894_/Q _06584_/C _06584_/D VGND VGND VPWR VPWR _06580_/X sky130_fd_sc_hd__and3_1
XFILLER_91_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14729_ _14746_/CLK _14729_/D VGND VGND VPWR VPWR _14729_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08250_ _08261_/A _08250_/B _08250_/C VGND VGND VPWR VPWR _08252_/B sky130_fd_sc_hd__and3_1
XFILLER_32_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07201_ _07201_/A VGND VGND VPWR VPWR _07205_/C sky130_fd_sc_hd__inv_2
X_08181_ _08167_/A _08170_/X _08180_/Y _07396_/A VGND VGND VPWR VPWR _08181_/X sky130_fd_sc_hd__a31o_1
XFILLER_119_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07132_ _07101_/A _07101_/B _07131_/Y VGND VGND VPWR VPWR _07133_/B sky130_fd_sc_hd__o21bai_1
X_07063_ _07063_/A _07063_/B _13707_/Q _07141_/C VGND VGND VPWR VPWR _07106_/A sky130_fd_sc_hd__and4_1
XFILLER_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06014_ _13583_/Q _13584_/Q _13585_/Q _13586_/Q VGND VGND VPWR VPWR _06017_/C sky130_fd_sc_hd__or4_1
XFILLER_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07965_ _07957_/A _07961_/X _07972_/C VGND VGND VPWR VPWR _07970_/B sky130_fd_sc_hd__a21oi_1
X_09704_ _09704_/A _09704_/B VGND VGND VPWR VPWR _09704_/X sky130_fd_sc_hd__and2_1
X_06916_ _07947_/B VGND VGND VPWR VPWR _06938_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_07896_ _07895_/B _07895_/C _13265_/Q VGND VGND VPWR VPWR _07904_/A sky130_fd_sc_hd__a21oi_1
XFILLER_110_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09635_ _09635_/A VGND VGND VPWR VPWR _12830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06847_ _06851_/A _06857_/A _06851_/B VGND VGND VPWR VPWR _06847_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_55_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09566_ _09574_/A _09574_/B _08733_/X VGND VGND VPWR VPWR _09566_/X sky130_fd_sc_hd__a21o_1
X_06778_ _06827_/A _06777_/B _06743_/A VGND VGND VPWR VPWR _06778_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08517_ _08642_/A VGND VGND VPWR VPWR _08517_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09497_ _13607_/Q _09525_/B VGND VGND VPWR VPWR _09498_/B sky130_fd_sc_hd__or2_1
XFILLER_12_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08448_ _13476_/Q VGND VGND VPWR VPWR _08544_/A sky130_fd_sc_hd__clkbuf_2
X_08379_ _08379_/A VGND VGND VPWR VPWR _12722_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10410_ _10410_/A _10410_/B VGND VGND VPWR VPWR _14217_/D sky130_fd_sc_hd__xnor2_1
XFILLER_149_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11390_ _13719_/Q _11394_/B VGND VGND VPWR VPWR _11391_/A sky130_fd_sc_hd__and2_1
XFILLER_164_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10341_ _13119_/D _10337_/B _10340_/A VGND VGND VPWR VPWR _10347_/A sky130_fd_sc_hd__a21oi_2
X_13060_ _13587_/CLK _13060_/D VGND VGND VPWR VPWR hold404/A sky130_fd_sc_hd__dfxtp_1
X_10272_ _10593_/A _14324_/Q VGND VGND VPWR VPWR _10272_/X sky130_fd_sc_hd__and2b_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12011_ _14313_/Q _12010_/X _12014_/S VGND VGND VPWR VPWR _12012_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13962_ _13972_/CLK _13962_/D VGND VGND VPWR VPWR _13962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12913_ _14737_/CLK _12913_/D VGND VGND VPWR VPWR _14695_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_73_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13893_ _14209_/CLK hold295/X VGND VGND VPWR VPWR _13893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _13799_/CLK _12844_/D VGND VGND VPWR VPWR hold335/A sky130_fd_sc_hd__dfxtp_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _13565_/CLK _12775_/D VGND VGND VPWR VPWR hold163/A sky130_fd_sc_hd__dfxtp_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _14608_/CLK _14514_/D VGND VGND VPWR VPWR _14514_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _11726_/A VGND VGND VPWR VPWR _14055_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14445_ _14598_/CLK _14445_/D VGND VGND VPWR VPWR _14445_/Q sky130_fd_sc_hd__dfxtp_1
X_11657_ _11691_/A VGND VGND VPWR VPWR _11708_/S sky130_fd_sc_hd__buf_2
X_10608_ _13964_/Q _13937_/Q _10607_/A VGND VGND VPWR VPWR _10608_/X sky130_fd_sc_hd__or3b_1
XFILLER_155_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14376_ _14536_/CLK _14377_/Q VGND VGND VPWR VPWR hold276/A sky130_fd_sc_hd__dfxtp_1
X_11588_ _11588_/A VGND VGND VPWR VPWR _13875_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13327_ _14709_/CLK _13327_/D VGND VGND VPWR VPWR _13327_/Q sky130_fd_sc_hd__dfxtp_4
X_10539_ _10539_/A _10539_/B VGND VGND VPWR VPWR _10539_/X sky130_fd_sc_hd__or2_1
XFILLER_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13258_ _13258_/CLK _13258_/D hold1/X VGND VGND VPWR VPWR _13258_/Q sky130_fd_sc_hd__dfrtp_4
X_12209_ _14120_/Q _14117_/Q _14121_/Q VGND VGND VPWR VPWR _12210_/C sky130_fd_sc_hd__a21o_1
X_13189_ _13606_/CLK _13189_/D VGND VGND VPWR VPWR hold405/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07750_ _07750_/A VGND VGND VPWR VPWR _07787_/B sky130_fd_sc_hd__inv_2
X_06701_ _07819_/B _06700_/Y _07909_/A VGND VGND VPWR VPWR _06702_/A sky130_fd_sc_hd__mux2_1
X_07681_ _07657_/A _07657_/B _07655_/B VGND VGND VPWR VPWR _07713_/B sky130_fd_sc_hd__a21oi_1
XFILLER_38_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09420_ _09420_/A _09420_/B _09420_/C _09420_/D VGND VGND VPWR VPWR _09421_/B sky130_fd_sc_hd__nor4_2
X_06632_ _13037_/Q VGND VGND VPWR VPWR _06704_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_25_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09351_ _09351_/A VGND VGND VPWR VPWR _12801_/D sky130_fd_sc_hd__clkbuf_1
X_06563_ _10337_/B _06563_/B _06563_/C VGND VGND VPWR VPWR _06565_/B sky130_fd_sc_hd__and3_1
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08302_ _08317_/C VGND VGND VPWR VPWR _08314_/B sky130_fd_sc_hd__clkbuf_1
X_09282_ _09282_/A _09282_/B _09276_/Y _09277_/X VGND VGND VPWR VPWR _09287_/C sky130_fd_sc_hd__or4bb_1
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06494_ _06488_/Y _06477_/B _06493_/Y VGND VGND VPWR VPWR _06499_/C sky130_fd_sc_hd__o21a_1
X_08233_ _08233_/A _08245_/A VGND VGND VPWR VPWR _08237_/A sky130_fd_sc_hd__or2_1
XFILLER_21_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08164_ _08164_/A _08164_/B _08164_/C VGND VGND VPWR VPWR _08166_/B sky130_fd_sc_hd__and3_1
XFILLER_20_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07115_ _07115_/A _07115_/B VGND VGND VPWR VPWR _07121_/A sky130_fd_sc_hd__xor2_1
XFILLER_118_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08095_ _12983_/Q _13283_/Q _08095_/S VGND VGND VPWR VPWR _08096_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07046_ _07031_/A _07163_/A _07044_/Y _07074_/A VGND VGND VPWR VPWR _07059_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08997_ _08997_/A _08997_/B VGND VGND VPWR VPWR _08997_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_29_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07948_ _07948_/A _07948_/B VGND VGND VPWR VPWR _07972_/A sky130_fd_sc_hd__nand2_1
XFILLER_29_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07879_ _07886_/C _07886_/D VGND VGND VPWR VPWR _07892_/D sky130_fd_sc_hd__or2_1
X_09618_ _13406_/Q _13604_/Q _09620_/S VGND VGND VPWR VPWR _09619_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10890_ _10890_/A VGND VGND VPWR VPWR _13203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09549_ _13615_/Q _09555_/B VGND VGND VPWR VPWR _09556_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12560_ _11370_/X _14725_/Q _12562_/S VGND VGND VPWR VPWR _12561_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11511_ _13838_/Q _11510_/X _11511_/S VGND VGND VPWR VPWR _11512_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12491_ _12491_/A VGND VGND VPWR VPWR _14675_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14230_ _14495_/CLK _14230_/D VGND VGND VPWR VPWR _14230_/Q sky130_fd_sc_hd__dfxtp_1
X_11442_ _13743_/Q _11444_/B VGND VGND VPWR VPWR _11443_/A sky130_fd_sc_hd__and2_1
XFILLER_109_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14161_ _14209_/CLK _14162_/Q VGND VGND VPWR VPWR _14161_/Q sky130_fd_sc_hd__dfxtp_1
X_11373_ _13844_/Q VGND VGND VPWR VPWR _11373_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13112_ _14634_/CLK _13112_/D VGND VGND VPWR VPWR _13112_/Q sky130_fd_sc_hd__dfxtp_1
X_10324_ _13747_/Q _13748_/Q VGND VGND VPWR VPWR _10330_/B sky130_fd_sc_hd__nor2_2
X_14092_ _14319_/CLK _14092_/D VGND VGND VPWR VPWR _14092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ _10190_/A _10242_/X _10246_/X VGND VGND VPWR VPWR _10255_/X sky130_fd_sc_hd__a21o_1
XFILLER_112_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13043_ _13525_/CLK _13043_/D VGND VGND VPWR VPWR _13076_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10186_ _10269_/S VGND VGND VPWR VPWR _14555_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_67_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13945_ _13945_/CLK _13945_/D VGND VGND VPWR VPWR _13945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13876_ _14656_/CLK _13876_/D VGND VGND VPWR VPWR _13876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12827_ _14327_/CLK _12827_/D VGND VGND VPWR VPWR hold251/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _13602_/CLK _12758_/D VGND VGND VPWR VPWR hold242/A sky130_fd_sc_hd__dfxtp_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11709_ _11709_/A VGND VGND VPWR VPWR _14036_/D sky130_fd_sc_hd__clkbuf_1
X_12689_ _13303_/CLK _12689_/D VGND VGND VPWR VPWR hold440/A sky130_fd_sc_hd__dfxtp_1
XFILLER_129_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14428_ _14644_/CLK _14428_/D VGND VGND VPWR VPWR _14428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14359_ _14536_/CLK _14359_/D VGND VGND VPWR VPWR _14359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08920_ _08889_/A _08889_/B _08919_/Y VGND VGND VPWR VPWR _08921_/B sky130_fd_sc_hd__o21bai_1
X_08851_ _08851_/A _08851_/B _13518_/D _08929_/C VGND VGND VPWR VPWR _08894_/A sky130_fd_sc_hd__and4_1
XFILLER_58_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07802_ _07802_/A _13252_/Q VGND VGND VPWR VPWR _07803_/B sky130_fd_sc_hd__nand2_1
X_05994_ _05994_/A _05994_/B VGND VGND VPWR VPWR _06231_/A sky130_fd_sc_hd__nor2_1
X_08782_ _08779_/Y _08780_/X _08775_/A _08776_/Y VGND VGND VPWR VPWR _08782_/X sky130_fd_sc_hd__a211o_1
X_07733_ _07733_/A _07733_/B VGND VGND VPWR VPWR _07734_/B sky130_fd_sc_hd__nand2_1
XFILLER_72_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07664_ _07664_/A _07664_/B VGND VGND VPWR VPWR _07708_/A sky130_fd_sc_hd__and2_1
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09403_ _09419_/C _09403_/B VGND VGND VPWR VPWR _09403_/X sky130_fd_sc_hd__xor2_1
X_06615_ _12904_/Q _06613_/A _06599_/X VGND VGND VPWR VPWR _06616_/B sky130_fd_sc_hd__o21ai_1
X_07595_ _13169_/D _07595_/B VGND VGND VPWR VPWR _11266_/B sky130_fd_sc_hd__xnor2_1
XFILLER_80_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09334_ _10831_/A VGND VGND VPWR VPWR _09343_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_80_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06546_ _12889_/Q _06552_/B VGND VGND VPWR VPWR _06547_/B sky130_fd_sc_hd__nor2_1
X_09265_ _09267_/B _09265_/B VGND VGND VPWR VPWR _09265_/Y sky130_fd_sc_hd__xnor2_1
X_06477_ _06488_/A _06477_/B VGND VGND VPWR VPWR _06477_/Y sky130_fd_sc_hd__xnor2_1
X_08216_ _08216_/A VGND VGND VPWR VPWR _13362_/D sky130_fd_sc_hd__clkbuf_1
X_09196_ _09195_/A _09220_/A _07524_/X VGND VGND VPWR VPWR _09196_/X sky130_fd_sc_hd__a21o_1
XFILLER_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08147_ _08147_/A _08147_/B VGND VGND VPWR VPWR _08147_/X sky130_fd_sc_hd__and2_1
XFILLER_106_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08078_ _12975_/Q _13275_/Q _08084_/S VGND VGND VPWR VPWR _08079_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07029_ _13112_/D VGND VGND VPWR VPWR _07086_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10040_ _13800_/Q _13784_/Q _13935_/D VGND VGND VPWR VPWR _10041_/A sky130_fd_sc_hd__mux2_1
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_130_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_103_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_29_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold65 hold65/A VGND VGND VPWR VPWR hold65/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_152_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold76 hold76/A VGND VGND VPWR VPWR hold76/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold87 hold87/A VGND VGND VPWR VPWR hold87/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_11991_ _14517_/Q VGND VGND VPWR VPWR _11991_/X sky130_fd_sc_hd__clkbuf_2
Xhold98 hold98/A VGND VGND VPWR VPWR hold98/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_56_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13730_ _13805_/CLK hold70/X VGND VGND VPWR VPWR _13730_/Q sky130_fd_sc_hd__dfxtp_1
X_10942_ _11092_/A VGND VGND VPWR VPWR _10942_/X sky130_fd_sc_hd__buf_2
XFILLER_45_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13661_ _13666_/CLK _13661_/D VGND VGND VPWR VPWR _13661_/Q sky130_fd_sc_hd__dfxtp_1
X_10873_ _10873_/A VGND VGND VPWR VPWR _13195_/D sky130_fd_sc_hd__clkbuf_1
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12612_ _14734_/Q _12611_/A _12633_/B VGND VGND VPWR VPWR _12612_/Y sky130_fd_sc_hd__a21boi_1
X_13592_ _13593_/CLK _13592_/D repeater56/X VGND VGND VPWR VPWR _13592_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_40_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12543_ _11326_/X _14717_/Q _12543_/S VGND VGND VPWR VPWR _12544_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12474_ _14668_/Q _12016_/A _12480_/S VGND VGND VPWR VPWR _12475_/A sky130_fd_sc_hd__mux2_1
X_14213_ _14440_/CLK _14213_/D VGND VGND VPWR VPWR _14213_/Q sky130_fd_sc_hd__dfxtp_1
X_11425_ _13735_/Q _11427_/B VGND VGND VPWR VPWR _11426_/A sky130_fd_sc_hd__and2_1
XANTENNA_7 input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14144_ _14159_/CLK _14197_/Q VGND VGND VPWR VPWR _14144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11356_ _11356_/A VGND VGND VPWR VPWR _13774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10307_ _10307_/A _10307_/B VGND VGND VPWR VPWR _13474_/D sky130_fd_sc_hd__nor2_1
XFILLER_3_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14075_ _14075_/CLK _14075_/D VGND VGND VPWR VPWR hold199/A sky130_fd_sc_hd__dfxtp_1
X_11287_ _11287_/A VGND VGND VPWR VPWR _13756_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ _14108_/CLK _13026_/D repeater59/X VGND VGND VPWR VPWR _13026_/Q sky130_fd_sc_hd__dfrtp_1
X_10238_ _14524_/D _10237_/X _14557_/D VGND VGND VPWR VPWR _10238_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10169_ _10160_/X _10168_/X _14293_/D VGND VGND VPWR VPWR _10169_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13928_ _14042_/CLK _13929_/Q VGND VGND VPWR VPWR _13928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13859_ _14656_/CLK _13859_/D VGND VGND VPWR VPWR _13859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06400_ _12910_/Q VGND VGND VPWR VPWR _06500_/A sky130_fd_sc_hd__clkinv_2
XFILLER_16_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07380_ _09139_/B _09139_/C _13140_/Q VGND VGND VPWR VPWR _07415_/A sky130_fd_sc_hd__a21oi_1
X_06331_ _14102_/Q _14086_/Q _06341_/S VGND VGND VPWR VPWR _06332_/A sky130_fd_sc_hd__mux2_1
X_09050_ _09050_/A VGND VGND VPWR VPWR _12760_/D sky130_fd_sc_hd__clkbuf_1
X_06262_ hold498/A _13974_/D VGND VGND VPWR VPWR _06262_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08001_ _13280_/Q _08001_/B VGND VGND VPWR VPWR _08003_/A sky130_fd_sc_hd__and2_1
XFILLER_116_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06193_ _06192_/X _06186_/X _06197_/A VGND VGND VPWR VPWR _06194_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold502 hold34/X VGND VGND VPWR VPWR hold502/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold513 hold14/X VGND VGND VPWR VPWR hold513/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09952_ _09952_/A VGND VGND VPWR VPWR _12862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08903_ _08903_/A _08903_/B VGND VGND VPWR VPWR _08909_/A sky130_fd_sc_hd__xor2_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _09885_/B _09883_/B _09883_/C VGND VGND VPWR VPWR _09884_/A sky130_fd_sc_hd__and3b_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08834_ _08819_/A _08951_/A _08832_/Y _08862_/A VGND VGND VPWR VPWR _08847_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08765_ _08706_/X _08767_/B _08763_/Y _08764_/X VGND VGND VPWR VPWR _13461_/D sky130_fd_sc_hd__a31o_1
X_05977_ _05977_/A _05977_/B _05977_/C VGND VGND VPWR VPWR _05977_/Y sky130_fd_sc_hd__nor3_1
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07716_ _07715_/B _07716_/B VGND VGND VPWR VPWR _07717_/B sky130_fd_sc_hd__and2b_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08696_ _09493_/A VGND VGND VPWR VPWR _08696_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07647_ _07701_/B _07668_/C _07723_/B _13244_/D VGND VGND VPWR VPWR _07649_/A sky130_fd_sc_hd__a22oi_1
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07578_ _07578_/A _07578_/B _07571_/Y _07572_/X VGND VGND VPWR VPWR _07583_/C sky130_fd_sc_hd__or4bb_1
XFILLER_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09317_ _13296_/Q _13534_/Q _09321_/S VGND VGND VPWR VPWR _09318_/A sky130_fd_sc_hd__mux2_1
X_06529_ _06529_/A _06529_/B VGND VGND VPWR VPWR _06529_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_21_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09248_ _09256_/A _09255_/A VGND VGND VPWR VPWR _09248_/X sky130_fd_sc_hd__or2_1
XFILLER_154_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_10_0_clk clkbuf_3_5_0_clk/X VGND VGND VPWR VPWR clkbuf_4_10_0_clk/X sky130_fd_sc_hd__clkbuf_2
X_09179_ _09189_/A _09180_/B VGND VGND VPWR VPWR _09186_/B sky130_fd_sc_hd__or2_1
XFILLER_5_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11210_ _14314_/Q _14484_/Q _14240_/Q _14070_/Q _11208_/X _11209_/X VGND VGND VPWR
+ VPWR _11210_/X sky130_fd_sc_hd__mux4_1
X_12190_ _14506_/Q _12007_/X _12194_/S VGND VGND VPWR VPWR _12191_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11141_ _11141_/A _11084_/X VGND VGND VPWR VPWR _11141_/X sky130_fd_sc_hd__or2b_1
Xoutput33 _13330_/Q VGND VGND VPWR VPWR data_o[12] sky130_fd_sc_hd__buf_2
XFILLER_123_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput44 _13340_/Q VGND VGND VPWR VPWR data_o[22] sky130_fd_sc_hd__buf_2
Xoutput55 _14729_/Q VGND VGND VPWR VPWR rts_o sky130_fd_sc_hd__buf_2
XFILLER_123_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11072_ _14605_/Q _14567_/Q _14498_/Q _14450_/Q _11044_/X _11045_/X VGND VGND VPWR
+ VPWR _11073_/A sky130_fd_sc_hd__mux4_1
XFILLER_49_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10023_ _10023_/A VGND VGND VPWR VPWR _10607_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11974_ _11974_/A VGND VGND VPWR VPWR _14301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13713_ _13727_/CLK hold45/X VGND VGND VPWR VPWR _13713_/Q sky130_fd_sc_hd__dfxtp_1
X_10925_ _11155_/A VGND VGND VPWR VPWR _10925_/X sky130_fd_sc_hd__clkbuf_1
X_14693_ _14693_/CLK _14693_/D VGND VGND VPWR VPWR _14693_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13644_ _14696_/CLK hold92/X VGND VGND VPWR VPWR _13644_/Q sky130_fd_sc_hd__dfxtp_1
X_10856_ _10856_/A VGND VGND VPWR VPWR _13187_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13575_ _14319_/CLK hold219/X VGND VGND VPWR VPWR _13575_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10787_ _10787_/A VGND VGND VPWR VPWR _13056_/D sky130_fd_sc_hd__clkbuf_1
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12526_ _11301_/X _14709_/Q _12532_/S VGND VGND VPWR VPWR _12527_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12457_ _14660_/Q _14517_/Q _12461_/S VGND VGND VPWR VPWR _12458_/A sky130_fd_sc_hd__mux2_1
X_11408_ _13727_/Q _11416_/B VGND VGND VPWR VPWR _11409_/A sky130_fd_sc_hd__and2_1
X_12388_ _14616_/Q _12016_/X _12394_/S VGND VGND VPWR VPWR _12389_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14127_ _14153_/CLK hold182/X VGND VGND VPWR VPWR hold429/A sky130_fd_sc_hd__dfxtp_1
XFILLER_113_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11339_ _11339_/A VGND VGND VPWR VPWR _13771_/D sky130_fd_sc_hd__clkbuf_1
X_14761__72 VGND VGND VPWR VPWR _14761__72/HI _13166_/D sky130_fd_sc_hd__conb_1
XFILLER_4_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14058_ _14495_/CLK _14058_/D VGND VGND VPWR VPWR _14058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05900_ _13811_/Q _13812_/Q _13813_/Q VGND VGND VPWR VPWR _05903_/A sky130_fd_sc_hd__or3_1
X_13009_ _13298_/CLK _13009_/D repeater59/X VGND VGND VPWR VPWR _13009_/Q sky130_fd_sc_hd__dfrtp_1
X_06880_ _06846_/B _06877_/Y _06878_/X _06879_/X VGND VGND VPWR VPWR _06899_/A sky130_fd_sc_hd__o211ai_4
XFILLER_67_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08550_ _08578_/A _08550_/B VGND VGND VPWR VPWR _08550_/X sky130_fd_sc_hd__or2_1
XFILLER_82_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07501_ _13151_/Q _07513_/B VGND VGND VPWR VPWR _07503_/A sky130_fd_sc_hd__nand2_1
XFILLER_35_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08481_ _08481_/A _08481_/B VGND VGND VPWR VPWR _08481_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_23_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07432_ _07438_/A _07442_/A VGND VGND VPWR VPWR _07434_/A sky130_fd_sc_hd__or2_1
XFILLER_62_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07363_ _07374_/A _07363_/B VGND VGND VPWR VPWR _07364_/B sky130_fd_sc_hd__and2_2
XFILLER_31_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09102_ _09095_/A _09095_/B _09101_/Y VGND VGND VPWR VPWR _09103_/B sky130_fd_sc_hd__o21ai_1
X_06314_ _06314_/A VGND VGND VPWR VPWR _14191_/D sky130_fd_sc_hd__clkbuf_1
X_07294_ _07294_/A _07294_/B VGND VGND VPWR VPWR _07294_/Y sky130_fd_sc_hd__xnor2_1
X_06245_ _14093_/Q _06245_/B VGND VGND VPWR VPWR _06246_/A sky130_fd_sc_hd__and2_1
X_09033_ _09033_/A VGND VGND VPWR VPWR _12752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06176_ _06176_/A VGND VGND VPWR VPWR _14175_/D sky130_fd_sc_hd__clkbuf_1
Xhold310 hold310/A VGND VGND VPWR VPWR hold310/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold321 hold321/A VGND VGND VPWR VPWR hold321/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold332 hold332/A VGND VGND VPWR VPWR hold332/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_117_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold343 hold343/A VGND VGND VPWR VPWR hold343/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold354 hold354/A VGND VGND VPWR VPWR hold354/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_105_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold365 hold365/A VGND VGND VPWR VPWR hold365/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold376 hold376/A VGND VGND VPWR VPWR hold376/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold387 hold387/A VGND VGND VPWR VPWR hold387/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold398 hold398/A VGND VGND VPWR VPWR hold398/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09935_ _13492_/Q _13681_/Q _09935_/S VGND VGND VPWR VPWR _09936_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ _13687_/Q _13688_/Q VGND VGND VPWR VPWR _09873_/D sky130_fd_sc_hd__and2_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ _13429_/Q VGND VGND VPWR VPWR _08874_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09797_ _13701_/Q VGND VGND VPWR VPWR _09834_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_85_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _08758_/A _08757_/A VGND VGND VPWR VPWR _08748_/Y sky130_fd_sc_hd__nand2_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _09550_/B VGND VGND VPWR VPWR _09562_/B sky130_fd_sc_hd__buf_2
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _10710_/A VGND VGND VPWR VPWR _12933_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11690_/A VGND VGND VPWR VPWR _14027_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10641_ _14194_/Q _14197_/Q VGND VGND VPWR VPWR _14145_/D sky130_fd_sc_hd__xor2_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13360_ _13434_/CLK _13360_/D repeater56/X VGND VGND VPWR VPWR _13360_/Q sky130_fd_sc_hd__dfrtp_1
X_10572_ _10572_/A VGND VGND VPWR VPWR _14438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12311_ _14571_/Q _11994_/X _12313_/S VGND VGND VPWR VPWR _12312_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13291_ _13296_/CLK hold352/X VGND VGND VPWR VPWR _13291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12242_ _11301_/X _14537_/Q _12248_/S VGND VGND VPWR VPWR _12243_/A sky130_fd_sc_hd__mux2_1
X_12173_ _12173_/A VGND VGND VPWR VPWR _14498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11124_ _13330_/Q _11079_/X _11113_/X _11123_/Y VGND VGND VPWR VPWR _13330_/D sky130_fd_sc_hd__o22a_1
XFILLER_111_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11055_ _14021_/Q _13987_/Q _13827_/Q _14539_/Q _11010_/X _11011_/X VGND VGND VPWR
+ VPWR _11056_/A sky130_fd_sc_hd__mux4_1
XFILLER_49_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10006_ _10006_/A VGND VGND VPWR VPWR _12669_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14745_ _14746_/CLK _14745_/D VGND VGND VPWR VPWR _14745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11957_ _14296_/Q _11956_/X _11966_/S VGND VGND VPWR VPWR _11958_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10908_ _14747_/Q VGND VGND VPWR VPWR _12590_/A sky130_fd_sc_hd__clkbuf_2
X_14676_ _14687_/CLK _14676_/D VGND VGND VPWR VPWR hold204/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11888_ _14241_/Q _11513_/X _11894_/S VGND VGND VPWR VPWR _11889_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13627_ _13635_/CLK hold381/X VGND VGND VPWR VPWR _13627_/Q sky130_fd_sc_hd__dfxtp_1
X_10839_ _13138_/Q _10841_/B VGND VGND VPWR VPWR _10840_/A sky130_fd_sc_hd__and2_1
X_13558_ _13558_/CLK hold151/X VGND VGND VPWR VPWR _13558_/Q sky130_fd_sc_hd__dfxtp_1
X_12509_ _12509_/A VGND VGND VPWR VPWR _14702_/D sky130_fd_sc_hd__clkbuf_1
X_13489_ _13722_/CLK hold315/X VGND VGND VPWR VPWR _13489_/Q sky130_fd_sc_hd__dfxtp_1
X_06030_ _14644_/Q _06030_/B VGND VGND VPWR VPWR _06361_/A sky130_fd_sc_hd__nand2_1
XFILLER_133_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07981_ _13277_/Q _07981_/B VGND VGND VPWR VPWR _07986_/B sky130_fd_sc_hd__xor2_1
XFILLER_141_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09720_ _09720_/A _09720_/B _09720_/C VGND VGND VPWR VPWR _09722_/B sky130_fd_sc_hd__and3_1
XFILLER_141_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06932_ _06932_/A _06932_/B VGND VGND VPWR VPWR _06936_/A sky130_fd_sc_hd__or2_1
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09651_ _13421_/Q _13619_/Q _09653_/S VGND VGND VPWR VPWR _09652_/A sky130_fd_sc_hd__mux2_1
X_06863_ _06863_/A _06863_/B VGND VGND VPWR VPWR _06863_/X sky130_fd_sc_hd__or2_1
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08602_ _08602_/A VGND VGND VPWR VPWR _09438_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_94_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09582_ _09577_/A _09578_/X _09581_/Y VGND VGND VPWR VPWR _09582_/Y sky130_fd_sc_hd__a21oi_1
X_06794_ _06794_/A _06794_/B _06827_/B VGND VGND VPWR VPWR _06794_/X sky130_fd_sc_hd__and3_1
X_08533_ _08517_/X _08531_/Y _08532_/X VGND VGND VPWR VPWR _13440_/D sky130_fd_sc_hd__o21bai_1
XFILLER_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08464_ _08633_/A VGND VGND VPWR VPWR _08464_/X sky130_fd_sc_hd__buf_2
XFILLER_50_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07415_ _07415_/A _07415_/B _07415_/C VGND VGND VPWR VPWR _07425_/C sky130_fd_sc_hd__or3_1
XFILLER_11_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08395_ _13094_/Q _13375_/Q _08395_/S VGND VGND VPWR VPWR _08396_/A sky130_fd_sc_hd__mux2_1
X_07346_ _13664_/Q _13660_/Q _13662_/Q _13658_/Q _13171_/Q _07344_/S VGND VGND VPWR
+ VPWR _07347_/B sky130_fd_sc_hd__mux4_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07277_ _07276_/B _07276_/C _07276_/A VGND VGND VPWR VPWR _07277_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09016_ _13209_/Q _13438_/Q _09018_/S VGND VGND VPWR VPWR _09017_/A sky130_fd_sc_hd__mux2_1
X_06228_ _06228_/A VGND VGND VPWR VPWR _14416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06159_ _14198_/D _14199_/D VGND VGND VPWR VPWR _06160_/A sky130_fd_sc_hd__or2_1
Xhold140 hold140/A VGND VGND VPWR VPWR hold140/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold151 hold151/A VGND VGND VPWR VPWR hold151/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold162 hold162/A VGND VGND VPWR VPWR hold162/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold173 hold173/A VGND VGND VPWR VPWR hold173/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold184 hold184/A VGND VGND VPWR VPWR hold184/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold195 hold195/A VGND VGND VPWR VPWR hold195/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09918_ _13484_/Q _13673_/Q _09924_/S VGND VGND VPWR VPWR _09919_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09849_ _13683_/Q _09851_/A _09848_/Y VGND VGND VPWR VPWR _13683_/D sky130_fd_sc_hd__o21a_1
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ _13805_/CLK _12860_/D VGND VGND VPWR VPWR hold341/A sky130_fd_sc_hd__dfxtp_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _13576_/Q _11817_/B VGND VGND VPWR VPWR _11812_/A sky130_fd_sc_hd__and2_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _13574_/CLK _12791_/D VGND VGND VPWR VPWR hold157/A sky130_fd_sc_hd__dfxtp_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14530_ _14530_/CLK hold132/X VGND VGND VPWR VPWR _14530_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _11742_/A VGND VGND VPWR VPWR _14062_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _14617_/CLK _14461_/D VGND VGND VPWR VPWR _14461_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11673_/A VGND VGND VPWR VPWR _14019_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13412_ _13617_/CLK hold443/X VGND VGND VPWR VPWR _13412_/Q sky130_fd_sc_hd__dfxtp_1
X_10624_ _14528_/Q _14363_/Q _14371_/Q hold17/X VGND VGND VPWR VPWR _10624_/X sky130_fd_sc_hd__or4_1
X_14392_ _14410_/CLK _14392_/D VGND VGND VPWR VPWR _14392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13343_ _14432_/CLK _13343_/D VGND VGND VPWR VPWR _13343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10555_ _10567_/A _10555_/B VGND VGND VPWR VPWR _10557_/C sky130_fd_sc_hd__and2_1
XFILLER_143_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13274_ _13274_/CLK _13274_/D repeater59/X VGND VGND VPWR VPWR _13274_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10486_ _10486_/A _10486_/B VGND VGND VPWR VPWR _10493_/A sky130_fd_sc_hd__or2_1
XFILLER_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12225_ _14126_/Q _12220_/X _12224_/Y VGND VGND VPWR VPWR _14519_/D sky130_fd_sc_hd__o21a_1
XFILLER_135_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12156_ _12156_/A VGND VGND VPWR VPWR _14490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11107_ _11088_/X _11104_/Y _11106_/Y _11095_/X VGND VGND VPWR VPWR _11108_/B sky130_fd_sc_hd__a211o_1
XFILLER_110_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12087_ _11359_/X _14461_/Q _12093_/S VGND VGND VPWR VPWR _12088_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11038_ _13324_/Q _11008_/X _11031_/X _11037_/Y VGND VGND VPWR VPWR _13324_/D sky130_fd_sc_hd__o22a_1
XFILLER_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12989_ _13351_/CLK _12989_/D VGND VGND VPWR VPWR hold515/A sky130_fd_sc_hd__dfxtp_2
X_14728_ _14737_/CLK _14728_/D VGND VGND VPWR VPWR _14728_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14659_ _14714_/CLK _14659_/D VGND VGND VPWR VPWR _14659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_180_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _14535_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_60_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07200_ _07200_/A VGND VGND VPWR VPWR _13350_/D sky130_fd_sc_hd__clkbuf_1
X_08180_ _13359_/Q _08180_/B VGND VGND VPWR VPWR _08180_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_158_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07131_ _07131_/A _07131_/B VGND VGND VPWR VPWR _07131_/Y sky130_fd_sc_hd__nor2_1
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07062_ _07063_/B _07165_/A _07190_/A _07063_/A VGND VGND VPWR VPWR _07064_/A sky130_fd_sc_hd__a22oi_1
XFILLER_145_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06013_ _13575_/Q _13580_/Q _13581_/Q _13582_/Q VGND VGND VPWR VPWR _06018_/C sky130_fd_sc_hd__or4_2
XFILLER_127_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07964_ _07970_/A _07964_/B VGND VGND VPWR VPWR _07972_/C sky130_fd_sc_hd__or2_1
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09703_ _14215_/Q _14213_/Q _09715_/S VGND VGND VPWR VPWR _09704_/B sky130_fd_sc_hd__mux2_1
X_06915_ _06861_/X _06919_/B _06914_/Y _06907_/X VGND VGND VPWR VPWR _13016_/D sky130_fd_sc_hd__a31o_1
XFILLER_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07895_ _13265_/Q _07895_/B _07895_/C VGND VGND VPWR VPWR _07905_/A sky130_fd_sc_hd__and3_1
X_09634_ _13413_/Q _13611_/Q _09642_/S VGND VGND VPWR VPWR _09635_/A sky130_fd_sc_hd__mux2_1
X_06846_ _06846_/A _06846_/B VGND VGND VPWR VPWR _06851_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09565_ _09574_/A _09574_/B VGND VGND VPWR VPWR _09565_/Y sky130_fd_sc_hd__nor2_1
X_06777_ _06827_/A _06777_/B VGND VGND VPWR VPWR _06794_/B sky130_fd_sc_hd__or2_1
X_08516_ _08504_/X _08530_/B _08513_/Y _08515_/X VGND VGND VPWR VPWR _13439_/D sky130_fd_sc_hd__a31o_1
X_09496_ _13607_/Q _09511_/B VGND VGND VPWR VPWR _09505_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08447_ _13475_/Q VGND VGND VPWR VPWR _08473_/C sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_171_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _14746_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08378_ _13086_/Q _13367_/Q _08384_/S VGND VGND VPWR VPWR _08379_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07329_ _07372_/S _13169_/Q VGND VGND VPWR VPWR _07329_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10340_ _10340_/A _10340_/B VGND VGND VPWR VPWR _13037_/D sky130_fd_sc_hd__nor2_1
X_10271_ _14595_/Q VGND VGND VPWR VPWR _10593_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12010_ _12010_/A VGND VGND VPWR VPWR _12010_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13961_ _13963_/CLK _13961_/D VGND VGND VPWR VPWR _13962_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_93_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12912_ _14536_/CLK _12912_/D VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13892_ _14209_/CLK hold95/X VGND VGND VPWR VPWR _13892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ _13721_/CLK _12843_/D VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _13704_/CLK _12774_/D VGND VGND VPWR VPWR hold268/A sky130_fd_sc_hd__dfxtp_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _14608_/CLK _14513_/D VGND VGND VPWR VPWR _14513_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11725_ _11294_/X _14055_/Q _11725_/S VGND VGND VPWR VPWR _11726_/A sky130_fd_sc_hd__mux2_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_162_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _14333_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14444_ _14652_/CLK _14444_/D VGND VGND VPWR VPWR _14444_/Q sky130_fd_sc_hd__dfxtp_1
X_11656_ _12226_/A _12342_/A VGND VGND VPWR VPWR _11691_/A sky130_fd_sc_hd__nor2_8
XFILLER_80_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10607_ _10607_/A _13945_/Q _13963_/Q VGND VGND VPWR VPWR _10607_/X sky130_fd_sc_hd__or3_1
X_14375_ _14536_/CLK hold276/X VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__dfxtp_1
X_11587_ _13651_/Q _11591_/B VGND VGND VPWR VPWR _11588_/A sky130_fd_sc_hd__and2_1
XFILLER_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13326_ _14657_/CLK _13326_/D VGND VGND VPWR VPWR _13326_/Q sky130_fd_sc_hd__dfxtp_4
X_10538_ _10539_/A _10539_/B VGND VGND VPWR VPWR _10540_/A sky130_fd_sc_hd__and2_1
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13257_ _13296_/CLK _13257_/D hold1/X VGND VGND VPWR VPWR _13257_/Q sky130_fd_sc_hd__dfrtp_2
X_10469_ _10469_/A _10468_/X VGND VGND VPWR VPWR _10471_/A sky130_fd_sc_hd__or2b_1
XFILLER_142_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12208_ _14120_/Q _14117_/Q _14121_/Q VGND VGND VPWR VPWR _12215_/C sky130_fd_sc_hd__and3_1
XFILLER_124_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13188_ _13423_/CLK _13188_/D VGND VGND VPWR VPWR hold453/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12139_ _14484_/Q _12013_/X _12139_/S VGND VGND VPWR VPWR _12140_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06700_ _06700_/A _06700_/B VGND VGND VPWR VPWR _06700_/Y sky130_fd_sc_hd__xnor2_1
X_07680_ _07680_/A _07680_/B VGND VGND VPWR VPWR _07713_/A sky130_fd_sc_hd__xnor2_1
XFILLER_37_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06631_ _13038_/Q VGND VGND VPWR VPWR _06671_/A sky130_fd_sc_hd__inv_2
XFILLER_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09350_ _13311_/Q _13549_/Q _09354_/S VGND VGND VPWR VPWR _09351_/A sky130_fd_sc_hd__mux2_1
X_06562_ _06562_/A VGND VGND VPWR VPWR _12890_/D sky130_fd_sc_hd__clkbuf_1
X_08301_ _13372_/Q _13373_/Q _08301_/C _08301_/D VGND VGND VPWR VPWR _08317_/C sky130_fd_sc_hd__and4_1
X_09281_ _13551_/Q _13552_/Q _07586_/B VGND VGND VPWR VPWR _09287_/B sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_153_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _14495_/CLK sky130_fd_sc_hd__clkbuf_16
X_06493_ _06493_/A _06493_/B VGND VGND VPWR VPWR _06493_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08232_ _13364_/Q _08232_/B VGND VGND VPWR VPWR _08245_/A sky130_fd_sc_hd__nor2_1
XFILLER_147_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08163_ _08161_/X _08114_/X _08162_/Y _08108_/X VGND VGND VPWR VPWR _08164_/C sky130_fd_sc_hd__o22a_1
XFILLER_119_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07114_ _07114_/A _07114_/B VGND VGND VPWR VPWR _07115_/B sky130_fd_sc_hd__or2_1
XFILLER_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08094_ _08094_/A VGND VGND VPWR VPWR _12706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07045_ _07119_/B _07141_/A _07045_/C VGND VGND VPWR VPWR _07074_/A sky130_fd_sc_hd__and3_1
XFILLER_133_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08996_ _08996_/A _08996_/B VGND VGND VPWR VPWR _08997_/B sky130_fd_sc_hd__xnor2_1
XFILLER_85_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07947_ _13272_/Q _07947_/B VGND VGND VPWR VPWR _07948_/B sky130_fd_sc_hd__or2_1
XFILLER_87_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07878_ _13263_/Q _07878_/B _07878_/C VGND VGND VPWR VPWR _07886_/D sky130_fd_sc_hd__and3_1
XFILLER_55_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09617_ _09617_/A VGND VGND VPWR VPWR _12822_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06829_ _06852_/A _06704_/X _06747_/Y VGND VGND VPWR VPWR _06829_/X sky130_fd_sc_hd__o21ba_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09548_ _09548_/A _09548_/B VGND VGND VPWR VPWR _09553_/C sky130_fd_sc_hd__nand2_1
XFILLER_24_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_144_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _14605_/CLK sky130_fd_sc_hd__clkbuf_16
X_09479_ _09460_/A _09466_/A _09467_/A VGND VGND VPWR VPWR _09479_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_24_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11510_ _12013_/A VGND VGND VPWR VPWR _11510_/X sky130_fd_sc_hd__clkbuf_2
X_12490_ _12496_/A _12496_/B hold499/X VGND VGND VPWR VPWR _12491_/A sky130_fd_sc_hd__and3_1
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11441_ _11441_/A VGND VGND VPWR VPWR _13811_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14160_ _14209_/CLK _14161_/Q VGND VGND VPWR VPWR _14160_/Q sky130_fd_sc_hd__dfxtp_1
X_11372_ _11372_/A VGND VGND VPWR VPWR _13777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13111_ _14634_/CLK hold515/X VGND VGND VPWR VPWR _13111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10323_ _13240_/D _13107_/Q _10322_/A VGND VGND VPWR VPWR _10329_/A sky130_fd_sc_hd__a21oi_1
X_14091_ _14098_/CLK _14091_/D VGND VGND VPWR VPWR _14091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13042_ _13525_/CLK _13042_/D VGND VGND VPWR VPWR _13075_/D sky130_fd_sc_hd__dfxtp_1
X_10254_ _10254_/A VGND VGND VPWR VPWR _14351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10185_ _10226_/A _14359_/Q VGND VGND VPWR VPWR _10269_/S sky130_fd_sc_hd__xor2_2
XFILLER_120_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13944_ _13964_/CLK _13944_/D VGND VGND VPWR VPWR _13944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13875_ _14656_/CLK _13875_/D VGND VGND VPWR VPWR _13875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12826_ _14327_/CLK _12826_/D VGND VGND VPWR VPWR hold149/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12757_ _13704_/CLK _12757_/D VGND VGND VPWR VPWR hold259/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_135_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _14050_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11708_ _14036_/Q _11522_/X _11708_/S VGND VGND VPWR VPWR _11709_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12688_ _13303_/CLK _12688_/D VGND VGND VPWR VPWR hold389/A sky130_fd_sc_hd__dfxtp_1
XFILLER_129_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14427_ _14536_/CLK _14427_/D VGND VGND VPWR VPWR _14427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11639_ _13995_/Q _11501_/X _11645_/S VGND VGND VPWR VPWR _11640_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14358_ _14425_/CLK _14358_/D VGND VGND VPWR VPWR _14358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13309_ _14275_/CLK hold74/X VGND VGND VPWR VPWR _13309_/Q sky130_fd_sc_hd__dfxtp_1
X_14289_ _14294_/CLK _14289_/D VGND VGND VPWR VPWR _14289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08850_ _08851_/B _08953_/A _08978_/A _08851_/A VGND VGND VPWR VPWR _08852_/A sky130_fd_sc_hd__a22oi_1
XFILLER_123_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07801_ _07801_/A VGND VGND VPWR VPWR _13666_/D sky130_fd_sc_hd__clkbuf_1
X_08781_ _08775_/A _08776_/Y _08779_/Y _08780_/X VGND VGND VPWR VPWR _08781_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_38_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05993_ _14096_/Q _14097_/Q _05993_/C _05993_/D VGND VGND VPWR VPWR _05994_/B sky130_fd_sc_hd__and4_1
XFILLER_97_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07732_ _07732_/A _07732_/B VGND VGND VPWR VPWR _07734_/A sky130_fd_sc_hd__xnor2_1
XFILLER_84_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07663_ _07663_/A VGND VGND VPWR VPWR _13658_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09402_ _09396_/A _09419_/A _09400_/Y _09401_/Y VGND VGND VPWR VPWR _09403_/B sky130_fd_sc_hd__a31o_1
X_06614_ _12903_/Q _12904_/Q _06620_/B VGND VGND VPWR VPWR _06616_/A sky130_fd_sc_hd__and3_1
XFILLER_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07594_ _07613_/A _07622_/A VGND VGND VPWR VPWR _07595_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09333_ _09333_/A VGND VGND VPWR VPWR _12793_/D sky130_fd_sc_hd__clkbuf_1
X_06545_ _12889_/Q _06552_/B VGND VGND VPWR VPWR _06547_/A sky130_fd_sc_hd__and2_1
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_126_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _13964_/CLK sky130_fd_sc_hd__clkbuf_16
X_09264_ _09264_/A _09264_/B VGND VGND VPWR VPWR _09265_/B sky130_fd_sc_hd__nand2_1
X_06476_ _06452_/A _06452_/B _06465_/A _06475_/Y VGND VGND VPWR VPWR _06477_/B sky130_fd_sc_hd__o31a_1
X_08215_ _08210_/B _08214_/Y _08215_/S VGND VGND VPWR VPWR _08216_/A sky130_fd_sc_hd__mux2_1
X_09195_ _09195_/A _09220_/A VGND VGND VPWR VPWR _09195_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08146_ _14007_/Q _14005_/Q _08161_/S VGND VGND VPWR VPWR _08147_/B sky130_fd_sc_hd__mux2_1
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08077_ _08077_/A VGND VGND VPWR VPWR _12698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07028_ _07028_/A _07028_/B VGND VGND VPWR VPWR _07032_/A sky130_fd_sc_hd__nor2_1
XFILLER_115_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_08979_ _08979_/A _08979_/B VGND VGND VPWR VPWR _08992_/B sky130_fd_sc_hd__nor2_1
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__clkbuf_1
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold66 hold66/A VGND VGND VPWR VPWR hold66/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold77 hold77/A VGND VGND VPWR VPWR hold77/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11990_ _11990_/A VGND VGND VPWR VPWR _14306_/D sky130_fd_sc_hd__clkbuf_1
Xhold88 hold88/A VGND VGND VPWR VPWR hold88/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_152_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold99 hold99/A VGND VGND VPWR VPWR hold99/X sky130_fd_sc_hd__buf_2
XFILLER_72_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10941_ _12584_/A VGND VGND VPWR VPWR _11092_/A sky130_fd_sc_hd__buf_4
XFILLER_90_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13660_ _13666_/CLK _13660_/D VGND VGND VPWR VPWR _13660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10872_ _13153_/Q _10874_/B VGND VGND VPWR VPWR _10873_/A sky130_fd_sc_hd__and2_1
XFILLER_71_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12611_ _12611_/A _12611_/B VGND VGND VPWR VPWR _14733_/D sky130_fd_sc_hd__nor2_1
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_117_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _13635_/CLK sky130_fd_sc_hd__clkbuf_16
X_13591_ _13593_/CLK _13591_/D repeater56/X VGND VGND VPWR VPWR _13591_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12542_ _12542_/A VGND VGND VPWR VPWR _14716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12473_ _12473_/A VGND VGND VPWR VPWR _14667_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14212_ _14212_/CLK _14212_/D VGND VGND VPWR VPWR _14212_/Q sky130_fd_sc_hd__dfxtp_1
X_11424_ _11424_/A VGND VGND VPWR VPWR _13803_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_8 input10/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14143_ _14294_/CLK _14143_/D VGND VGND VPWR VPWR _14143_/Q sky130_fd_sc_hd__dfxtp_1
X_11355_ _13774_/Q _11354_/X _11355_/S VGND VGND VPWR VPWR _11356_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10306_ _10306_/A _13511_/D _10306_/C VGND VGND VPWR VPWR _10307_/B sky130_fd_sc_hd__nor3_1
XFILLER_153_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14074_ _14726_/CLK _14074_/D VGND VGND VPWR VPWR _14074_/Q sky130_fd_sc_hd__dfxtp_1
X_11286_ _13756_/Q _11285_/X _11295_/S VGND VGND VPWR VPWR _11287_/A sky130_fd_sc_hd__mux2_1
X_13025_ _13027_/CLK _13025_/D repeater59/X VGND VGND VPWR VPWR _13025_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10237_ _10237_/A _10237_/B VGND VGND VPWR VPWR _10237_/X sky130_fd_sc_hd__or2_1
XFILLER_79_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10168_ _10103_/A _10155_/X _10159_/X VGND VGND VPWR VPWR _10168_/X sky130_fd_sc_hd__a21o_1
XFILLER_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10099_ _10182_/S VGND VGND VPWR VPWR _14292_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_75_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13927_ _14042_/CLK _13928_/Q VGND VGND VPWR VPWR hold93/A sky130_fd_sc_hd__dfxtp_1
XFILLER_81_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13858_ _14180_/CLK _13858_/D VGND VGND VPWR VPWR _13858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12809_ _13635_/CLK _12809_/D VGND VGND VPWR VPWR hold387/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_108_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _13604_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13789_ _13799_/CLK _13789_/D VGND VGND VPWR VPWR _13789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06330_ _06330_/A VGND VGND VPWR VPWR _14426_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06261_ _06259_/A _06259_/Y _13965_/D _06260_/X VGND VGND VPWR VPWR _13975_/D sky130_fd_sc_hd__a22o_1
XFILLER_129_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08000_ _07987_/A _07987_/B _07998_/Y _07999_/X VGND VGND VPWR VPWR _08013_/A sky130_fd_sc_hd__a31oi_2
X_06192_ _14419_/Q _14417_/Q _14426_/Q VGND VGND VPWR VPWR _06192_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold503 hold503/A VGND VGND VPWR VPWR hold503/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold514 hold514/A VGND VGND VPWR VPWR hold514/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_116_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09951_ _13499_/Q _13688_/Q _09957_/S VGND VGND VPWR VPWR _09952_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08902_ _08902_/A _08902_/B VGND VGND VPWR VPWR _08903_/B sky130_fd_sc_hd__or2_1
XFILLER_143_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _13691_/Q _13692_/Q _09881_/D _13693_/Q VGND VGND VPWR VPWR _09883_/C sky130_fd_sc_hd__a31o_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08833_ _08907_/B _08929_/A _08833_/C VGND VGND VPWR VPWR _08862_/A sky130_fd_sc_hd__and3_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08764_ _09506_/A VGND VGND VPWR VPWR _08764_/X sky130_fd_sc_hd__buf_2
X_05976_ _05976_/A _05976_/B _05976_/C VGND VGND VPWR VPWR _05977_/C sky130_fd_sc_hd__or3_1
XFILLER_54_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07715_ _07716_/B _07715_/B VGND VGND VPWR VPWR _07735_/B sky130_fd_sc_hd__and2b_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08695_ _08698_/A _08714_/B VGND VGND VPWR VPWR _08695_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07646_ _07646_/A _07688_/A VGND VGND VPWR VPWR _07664_/A sky130_fd_sc_hd__nor2_1
XFILLER_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07577_ _13159_/Q _13160_/Q _07586_/B VGND VGND VPWR VPWR _07583_/B sky130_fd_sc_hd__o21ai_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09316_ _09316_/A VGND VGND VPWR VPWR _12785_/D sky130_fd_sc_hd__clkbuf_1
X_06528_ _06527_/Y _06520_/B _06515_/A VGND VGND VPWR VPWR _06529_/B sky130_fd_sc_hd__a21oi_1
X_09247_ _09256_/A _09255_/A VGND VGND VPWR VPWR _09247_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06459_ _06443_/X _06458_/X _06395_/X _06444_/Y VGND VGND VPWR VPWR _06460_/C sky130_fd_sc_hd__o22a_1
XFILLER_31_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09178_ _09173_/A _09173_/B _09177_/X _09172_/B VGND VGND VPWR VPWR _09180_/B sky130_fd_sc_hd__a31o_1
XFILLER_147_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08129_ _14006_/Q _14004_/Q _13424_/Q VGND VGND VPWR VPWR _08129_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11140_ _14027_/Q _13993_/Q _13833_/Q _14545_/Q _11081_/X _11082_/X VGND VGND VPWR
+ VPWR _11141_/A sky130_fd_sc_hd__mux4_1
XFILLER_122_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput34 _13331_/Q VGND VGND VPWR VPWR data_o[13] sky130_fd_sc_hd__buf_2
XFILLER_123_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput45 _13341_/Q VGND VGND VPWR VPWR data_o[23] sky130_fd_sc_hd__buf_2
XFILLER_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11071_ _11065_/X _11068_/X _11070_/X _11015_/X VGND VGND VPWR VPWR _11071_/X sky130_fd_sc_hd__o211a_1
XFILLER_122_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10022_ _13948_/Q _13940_/Q _10023_/A VGND VGND VPWR VPWR _10606_/C sky130_fd_sc_hd__mux2_1
XFILLER_76_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11973_ _14301_/Q _11972_/X _11982_/S VGND VGND VPWR VPWR _11974_/A sky130_fd_sc_hd__mux2_1
X_10924_ _12590_/A VGND VGND VPWR VPWR _11155_/A sky130_fd_sc_hd__clkbuf_4
X_13712_ _14256_/CLK _13712_/D VGND VGND VPWR VPWR _13712_/Q sky130_fd_sc_hd__dfxtp_1
X_14692_ _14692_/CLK hold191/X VGND VGND VPWR VPWR hold280/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13643_ _13653_/CLK hold445/X VGND VGND VPWR VPWR _13643_/Q sky130_fd_sc_hd__dfxtp_1
X_10855_ _13145_/Q _10863_/B VGND VGND VPWR VPWR _10856_/A sky130_fd_sc_hd__and2_1
XFILLER_32_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13574_ _13574_/CLK hold269/X VGND VGND VPWR VPWR _13574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10786_ _13014_/Q _10790_/B VGND VGND VPWR VPWR _10787_/A sky130_fd_sc_hd__and2_1
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12525_ _12525_/A VGND VGND VPWR VPWR _14708_/D sky130_fd_sc_hd__clkbuf_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12456_ _12456_/A VGND VGND VPWR VPWR _14659_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11407_ _11429_/A VGND VGND VPWR VPWR _11416_/B sky130_fd_sc_hd__clkbuf_1
X_12387_ _12387_/A VGND VGND VPWR VPWR _14615_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14126_ _14292_/CLK hold243/X VGND VGND VPWR VPWR _14126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11338_ _13771_/Q _11337_/X _11355_/S VGND VGND VPWR VPWR _11339_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14057_ _14600_/CLK _14057_/D VGND VGND VPWR VPWR _14057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11269_ _11269_/A VGND VGND VPWR VPWR _13712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13008_ _13264_/CLK _13008_/D repeater59/X VGND VGND VPWR VPWR _13008_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07500_ _07495_/X _07497_/X _07498_/Y _07499_/X VGND VGND VPWR VPWR _13150_/D sky130_fd_sc_hd__a31o_1
X_08480_ _08477_/Y _08480_/B VGND VGND VPWR VPWR _08481_/B sky130_fd_sc_hd__and2b_1
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07431_ _07435_/A _07435_/B _13144_/Q VGND VGND VPWR VPWR _07442_/A sky130_fd_sc_hd__a21oi_1
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07362_ _07327_/X _07224_/A _07241_/A VGND VGND VPWR VPWR _07363_/B sky130_fd_sc_hd__o21a_1
XFILLER_149_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09101_ _13525_/Q _09101_/B VGND VGND VPWR VPWR _09101_/Y sky130_fd_sc_hd__nand2_1
X_06313_ _13877_/Q _13861_/Q _06313_/S VGND VGND VPWR VPWR _06314_/A sky130_fd_sc_hd__mux2_1
X_07293_ _07276_/A _07276_/B _07292_/Y VGND VGND VPWR VPWR _07294_/B sky130_fd_sc_hd__o21ai_1
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09032_ _13216_/Q _13445_/Q _09040_/S VGND VGND VPWR VPWR _09033_/A sky130_fd_sc_hd__mux2_1
X_06244_ _06244_/A VGND VGND VPWR VPWR _14391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold300 hold300/A VGND VGND VPWR VPWR hold300/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06175_ _13861_/Q _06175_/B VGND VGND VPWR VPWR _06176_/A sky130_fd_sc_hd__and2_1
Xhold311 hold311/A VGND VGND VPWR VPWR hold311/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold322 hold322/A VGND VGND VPWR VPWR hold322/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold333 hold333/A VGND VGND VPWR VPWR hold333/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_105_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold344 hold344/A VGND VGND VPWR VPWR hold344/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold355 hold355/A VGND VGND VPWR VPWR hold355/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_117_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold366 hold366/A VGND VGND VPWR VPWR hold366/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold377 hold377/A VGND VGND VPWR VPWR hold377/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold388 hold388/A VGND VGND VPWR VPWR hold388/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09934_ _09934_/A VGND VGND VPWR VPWR _12854_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold399 hold399/A VGND VGND VPWR VPWR hold399/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_113_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09865_ _09865_/A _09865_/B VGND VGND VPWR VPWR _13687_/D sky130_fd_sc_hd__nor2_1
XFILLER_98_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ _08816_/A _08816_/B VGND VGND VPWR VPWR _08820_/A sky130_fd_sc_hd__nor2_1
XFILLER_46_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09796_ _09796_/A _09796_/B VGND VGND VPWR VPWR _09796_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_86_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08747_ _13459_/Q _09542_/B VGND VGND VPWR VPWR _08757_/A sky130_fd_sc_hd__xor2_1
XFILLER_27_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05959_ _13643_/Q _13644_/Q _13645_/Q _05959_/D VGND VGND VPWR VPWR _05959_/X sky130_fd_sc_hd__and4_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08678_ _08746_/A VGND VGND VPWR VPWR _09550_/B sky130_fd_sc_hd__buf_2
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07629_ _07626_/Y _07656_/A _14702_/Q _07745_/A VGND VGND VPWR VPWR _07656_/B sky130_fd_sc_hd__and4bb_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10640_ _13933_/Q _10640_/B VGND VGND VPWR VPWR _13909_/D sky130_fd_sc_hd__xnor2_1
XFILLER_22_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10571_ _10575_/B _10571_/B VGND VGND VPWR VPWR _10572_/A sky130_fd_sc_hd__and2_1
XFILLER_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12310_ _12310_/A VGND VGND VPWR VPWR _14570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13290_ _13296_/CLK hold382/X VGND VGND VPWR VPWR _13290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12241_ _12241_/A VGND VGND VPWR VPWR _14536_/D sky130_fd_sc_hd__clkbuf_1
X_12172_ _14498_/Q _11981_/X _12172_/S VGND VGND VPWR VPWR _12173_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11123_ _11179_/A _11123_/B VGND VGND VPWR VPWR _11123_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11054_ _14303_/Q _14473_/Q _14229_/Q _14059_/Q _10993_/X _10995_/X VGND VGND VPWR
+ VPWR _11054_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10005_ _10004_/X _10001_/X _10635_/B VGND VGND VPWR VPWR _10006_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14744_ _14749_/CLK _14744_/D VGND VGND VPWR VPWR _14744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11956_ _14695_/Q VGND VGND VPWR VPWR _11956_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10907_ _12626_/B VGND VGND VPWR VPWR _10907_/X sky130_fd_sc_hd__clkbuf_2
X_14675_ _14688_/CLK _14675_/D VGND VGND VPWR VPWR hold345/A sky130_fd_sc_hd__dfxtp_1
X_11887_ _11887_/A VGND VGND VPWR VPWR _14240_/D sky130_fd_sc_hd__clkbuf_1
X_13626_ _13626_/CLK hold128/X VGND VGND VPWR VPWR _13626_/Q sky130_fd_sc_hd__dfxtp_1
X_10838_ _10838_/A VGND VGND VPWR VPWR _13179_/D sky130_fd_sc_hd__clkbuf_1
X_13557_ _13558_/CLK hold174/X VGND VGND VPWR VPWR _13557_/Q sky130_fd_sc_hd__dfxtp_1
X_10769_ _10769_/A VGND VGND VPWR VPWR _13048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12508_ _10592_/B _12508_/B VGND VGND VPWR VPWR _12509_/A sky130_fd_sc_hd__and2b_1
X_13488_ _13722_/CLK hold35/X VGND VGND VPWR VPWR _13488_/Q sky130_fd_sc_hd__dfxtp_1
X_12439_ _14652_/Q _14698_/Q _12439_/S VGND VGND VPWR VPWR _12440_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14109_ _14319_/CLK _14109_/D VGND VGND VPWR VPWR _14109_/Q sky130_fd_sc_hd__dfxtp_1
X_07980_ _07978_/Y _07979_/X _07932_/X VGND VGND VPWR VPWR _13276_/D sky130_fd_sc_hd__a21o_1
X_06931_ _06932_/B _06929_/X _06930_/X VGND VGND VPWR VPWR _13018_/D sky130_fd_sc_hd__o21bai_1
XFILLER_68_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09650_ _09650_/A VGND VGND VPWR VPWR _12837_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06862_ _13012_/Q _07902_/B VGND VGND VPWR VPWR _06870_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08601_ _08620_/A _08601_/B VGND VGND VPWR VPWR _08601_/X sky130_fd_sc_hd__xor2_1
X_09581_ _13620_/Q _09581_/B VGND VGND VPWR VPWR _09581_/Y sky130_fd_sc_hd__xnor2_1
X_06793_ _06793_/A _06793_/B VGND VGND VPWR VPWR _06793_/Y sky130_fd_sc_hd__nand2_1
X_08532_ _08733_/A _08532_/B _08536_/A VGND VGND VPWR VPWR _08532_/X sky130_fd_sc_hd__and3_1
XFILLER_24_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08463_ _09422_/S VGND VGND VPWR VPWR _08633_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07414_ _07414_/A _07414_/B _07414_/C VGND VGND VPWR VPWR _07415_/C sky130_fd_sc_hd__or3_1
XFILLER_149_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08394_ _08394_/A VGND VGND VPWR VPWR _12729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07345_ _07428_/A _07344_/X _07329_/Y VGND VGND VPWR VPWR _07345_/X sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_30_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _13303_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_136_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07276_ _07276_/A _07276_/B _07276_/C VGND VGND VPWR VPWR _07276_/X sky130_fd_sc_hd__or3_1
XFILLER_136_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09015_ _09015_/A VGND VGND VPWR VPWR _12744_/D sky130_fd_sc_hd__clkbuf_1
X_06227_ _10626_/B _06226_/X _10208_/S VGND VGND VPWR VPWR _06228_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold130 hold130/A VGND VGND VPWR VPWR hold130/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06158_ _06158_/A VGND VGND VPWR VPWR _14199_/D sky130_fd_sc_hd__clkbuf_1
Xhold141 hold141/A VGND VGND VPWR VPWR hold141/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold152 hold152/A VGND VGND VPWR VPWR hold152/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold163 hold163/A VGND VGND VPWR VPWR hold163/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold174 hold174/A VGND VGND VPWR VPWR hold174/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold185 hold185/A VGND VGND VPWR VPWR hold185/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06089_ _13966_/D _13967_/D VGND VGND VPWR VPWR _06090_/A sky130_fd_sc_hd__or2_1
Xhold196 hold196/A VGND VGND VPWR VPWR hold196/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09917_ _09917_/A VGND VGND VPWR VPWR _12846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_97_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _13680_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ _13683_/Q _09851_/A _09672_/Y VGND VGND VPWR VPWR _09848_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _13676_/Q _09785_/B VGND VGND VPWR VPWR _09793_/A sky130_fd_sc_hd__nor2_1
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _11810_/A VGND VGND VPWR VPWR _14097_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _13570_/CLK _12790_/D VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__dfxtp_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11741_ _11317_/X _14062_/Q _11747_/S VGND VGND VPWR VPWR _11742_/A sky130_fd_sc_hd__mux2_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _14019_/Q _11469_/X _11678_/S VGND VGND VPWR VPWR _11673_/A sky130_fd_sc_hd__mux2_1
X_14460_ _14579_/CLK _14460_/D VGND VGND VPWR VPWR _14460_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10623_ _14520_/Q _14530_/Q VGND VGND VPWR VPWR _10623_/X sky130_fd_sc_hd__and2_1
X_13411_ _13617_/CLK hold424/X VGND VGND VPWR VPWR _13411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14391_ _14732_/CLK _14391_/D VGND VGND VPWR VPWR _14391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_21_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _13552_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13342_ _14432_/CLK _13342_/D VGND VGND VPWR VPWR _13342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10554_ _10557_/B VGND VGND VPWR VPWR _10573_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13273_ _13273_/CLK _13273_/D repeater59/X VGND VGND VPWR VPWR _13273_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10485_ _10485_/A _10485_/B _10485_/C VGND VGND VPWR VPWR _10486_/B sky130_fd_sc_hd__and3_1
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12224_ _14126_/Q _12220_/X _12205_/X VGND VGND VPWR VPWR _12224_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_108_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12155_ _14490_/Q _11956_/X _12161_/S VGND VGND VPWR VPWR _12156_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11106_ _11106_/A _11106_/B VGND VGND VPWR VPWR _11106_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12086_ _12086_/A VGND VGND VPWR VPWR _14460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_88_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _14440_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11037_ _11037_/A _11037_/B VGND VGND VPWR VPWR _11037_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12988_ _14636_/CLK _12988_/D VGND VGND VPWR VPWR _13109_/D sky130_fd_sc_hd__dfxtp_2
X_14727_ _14746_/CLK _14727_/D VGND VGND VPWR VPWR _14727_/Q sky130_fd_sc_hd__dfxtp_1
X_11939_ _11939_/A VGND VGND VPWR VPWR _14275_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14658_ _14714_/CLK _14658_/D VGND VGND VPWR VPWR _14658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13609_ _13610_/CLK _13609_/D repeater57/X VGND VGND VPWR VPWR _13609_/Q sky130_fd_sc_hd__dfrtp_2
X_14589_ _14678_/CLK _14687_/Q VGND VGND VPWR VPWR _14589_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_12_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _13570_/CLK sky130_fd_sc_hd__clkbuf_16
X_07130_ _07153_/A _07130_/B VGND VGND VPWR VPWR _07134_/B sky130_fd_sc_hd__or2_1
XFILLER_9_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07061_ _07141_/C VGND VGND VPWR VPWR _07190_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06012_ _06012_/A _06012_/B _06012_/C VGND VGND VPWR VPWR _06012_/X sky130_fd_sc_hd__and3_1
XFILLER_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07963_ _13274_/Q _07963_/B VGND VGND VPWR VPWR _07964_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_79_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _14688_/CLK sky130_fd_sc_hd__clkbuf_16
X_06914_ _06914_/A _06914_/B _06924_/C VGND VGND VPWR VPWR _06914_/Y sky130_fd_sc_hd__nand3_1
X_09702_ _09787_/S _09700_/X _09701_/X _09767_/A VGND VGND VPWR VPWR _09702_/X sky130_fd_sc_hd__o211a_1
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07894_ _07811_/X _07898_/B _07893_/Y _06838_/X VGND VGND VPWR VPWR _13264_/D sky130_fd_sc_hd__a31o_1
XFILLER_114_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09633_ _09644_/A VGND VGND VPWR VPWR _09642_/S sky130_fd_sc_hd__clkbuf_2
X_06845_ _06840_/A _06843_/A _13011_/Q VGND VGND VPWR VPWR _06857_/A sky130_fd_sc_hd__a21oi_1
XFILLER_82_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09564_ _09564_/A _09564_/B VGND VGND VPWR VPWR _09574_/B sky130_fd_sc_hd__or2_1
X_06776_ _06740_/X _06775_/Y _06759_/A VGND VGND VPWR VPWR _06777_/B sky130_fd_sc_hd__a21o_1
XFILLER_36_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08515_ _08665_/A _09394_/B VGND VGND VPWR VPWR _08515_/X sky130_fd_sc_hd__and2_1
XFILLER_36_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09495_ _09495_/A _09491_/B VGND VGND VPWR VPWR _09500_/B sky130_fd_sc_hd__or2b_1
XFILLER_70_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08446_ _08506_/S _13712_/Q VGND VGND VPWR VPWR _08446_/X sky130_fd_sc_hd__and2b_1
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08377_ _08377_/A VGND VGND VPWR VPWR _12721_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07328_ _13169_/Q _13665_/Q _07344_/S VGND VGND VPWR VPWR _07328_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07259_ _13165_/Q VGND VGND VPWR VPWR _07473_/A sky130_fd_sc_hd__inv_2
XFILLER_137_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10270_ _10270_/A VGND VGND VPWR VPWR _14356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13960_ _14196_/CLK _13960_/D VGND VGND VPWR VPWR hold156/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12911_ _12970_/CLK _12911_/D VGND VGND VPWR VPWR _12911_/Q sky130_fd_sc_hd__dfxtp_1
X_13891_ _14693_/CLK hold339/X VGND VGND VPWR VPWR _13891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _13727_/CLK _12842_/D VGND VGND VPWR VPWR hold414/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _13626_/CLK _12773_/D VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__dfxtp_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14615_/CLK _14512_/D VGND VGND VPWR VPWR _14512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _11724_/A VGND VGND VPWR VPWR _14054_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _11655_/A _11712_/B _12582_/A VGND VGND VPWR VPWR _12342_/A sky130_fd_sc_hd__or3_4
X_14443_ _14598_/CLK _14443_/D VGND VGND VPWR VPWR _14443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10606_ _10606_/A _10606_/B _10606_/C _10606_/D VGND VGND VPWR VPWR _10606_/X sky130_fd_sc_hd__or4_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11586_ _11586_/A VGND VGND VPWR VPWR _13874_/D sky130_fd_sc_hd__clkbuf_1
X_14374_ _14710_/CLK hold20/X VGND VGND VPWR VPWR _14374_/Q sky130_fd_sc_hd__dfxtp_1
X_10537_ _10537_/A _10537_/B VGND VGND VPWR VPWR _10539_/B sky130_fd_sc_hd__xnor2_1
X_13325_ _14657_/CLK _13325_/D VGND VGND VPWR VPWR _13325_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_7_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10468_ _10468_/A _10468_/B VGND VGND VPWR VPWR _10468_/X sky130_fd_sc_hd__or2_1
X_13256_ _13256_/CLK _13256_/D hold1/X VGND VGND VPWR VPWR _13256_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12207_ _14120_/Q _14117_/Q _12206_/Y VGND VGND VPWR VPWR _14513_/D sky130_fd_sc_hd__a21oi_1
X_13187_ _13423_/CLK _13187_/D VGND VGND VPWR VPWR hold348/A sky130_fd_sc_hd__dfxtp_1
X_10399_ _10415_/A _10376_/A _10374_/A _10411_/B VGND VGND VPWR VPWR _10400_/B sky130_fd_sc_hd__a31o_1
X_12138_ _12138_/A VGND VGND VPWR VPWR _14483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12069_ _12069_/A VGND VGND VPWR VPWR _14452_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_1_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _14722_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06630_ _06630_/A VGND VGND VPWR VPWR _06881_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_25_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06561_ _06556_/B _06560_/Y _06599_/A VGND VGND VPWR VPWR _06562_/A sky130_fd_sc_hd__mux2_1
X_08300_ _13372_/Q _08294_/X _08299_/Y VGND VGND VPWR VPWR _13372_/D sky130_fd_sc_hd__a21oi_1
XFILLER_33_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09280_ _08218_/X _09278_/Y _09279_/X _09215_/X VGND VGND VPWR VPWR _13552_/D sky130_fd_sc_hd__a31o_1
X_06492_ _06492_/A VGND VGND VPWR VPWR _12883_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08231_ _13364_/Q _08231_/B _08279_/D VGND VGND VPWR VPWR _08233_/A sky130_fd_sc_hd__and3_1
X_08162_ _08176_/A _08162_/B VGND VGND VPWR VPWR _08162_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07113_ _07113_/A _07113_/B VGND VGND VPWR VPWR _07115_/A sky130_fd_sc_hd__xnor2_1
X_08093_ _12982_/Q _13282_/Q _08095_/S VGND VGND VPWR VPWR _08094_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07044_ _07063_/B _07119_/B _07141_/A _07119_/A VGND VGND VPWR VPWR _07044_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08995_ _08995_/A _08995_/B VGND VGND VPWR VPWR _08996_/B sky130_fd_sc_hd__xnor2_1
XFILLER_75_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07946_ _13272_/Q _07955_/B VGND VGND VPWR VPWR _07948_/A sky130_fd_sc_hd__nand2_1
XFILLER_130_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07877_ _07878_/B _07878_/C _13263_/Q VGND VGND VPWR VPWR _07886_/C sky130_fd_sc_hd__a21oi_1
XFILLER_141_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09616_ _13405_/Q _13603_/Q _09620_/S VGND VGND VPWR VPWR _09617_/A sky130_fd_sc_hd__mux2_1
X_06828_ _06740_/X _06775_/Y _06826_/C _06827_/X _06759_/A VGND VGND VPWR VPWR _06828_/X
+ sky130_fd_sc_hd__a2111o_1
X_09547_ _09547_/A _09547_/B VGND VGND VPWR VPWR _09548_/B sky130_fd_sc_hd__and2_1
X_06759_ _06759_/A _06775_/B VGND VGND VPWR VPWR _06762_/A sky130_fd_sc_hd__or2_1
X_09478_ _09478_/A _09478_/B VGND VGND VPWR VPWR _09478_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08429_ _13474_/Q VGND VGND VPWR VPWR _08506_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_8_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11440_ _13742_/Q _11444_/B VGND VGND VPWR VPWR _11441_/A sky130_fd_sc_hd__and2_1
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11371_ _13777_/Q _11370_/X _11376_/S VGND VGND VPWR VPWR _11372_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13110_ _14645_/CLK hold187/X VGND VGND VPWR VPWR _13110_/Q sky130_fd_sc_hd__dfxtp_1
X_10322_ _10322_/A _10322_/B VGND VGND VPWR VPWR _13170_/D sky130_fd_sc_hd__nor2_1
XFILLER_164_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14090_ _14098_/CLK _14090_/D VGND VGND VPWR VPWR _14090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13041_ _14636_/CLK _13041_/D VGND VGND VPWR VPWR hold494/A sky130_fd_sc_hd__dfxtp_1
X_10253_ _10248_/X _10252_/X _14555_/D VGND VGND VPWR VPWR _10254_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10184_ _14358_/Q VGND VGND VPWR VPWR _10226_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_132_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13943_ _13963_/CLK _13943_/D VGND VGND VPWR VPWR _13943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13874_ _14656_/CLK _13874_/D VGND VGND VPWR VPWR _13874_/Q sky130_fd_sc_hd__dfxtp_1
X_12825_ _14327_/CLK _12825_/D VGND VGND VPWR VPWR hold407/A sky130_fd_sc_hd__dfxtp_1
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _13722_/CLK _12756_/D VGND VGND VPWR VPWR hold218/A sky130_fd_sc_hd__dfxtp_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11707_ _11707_/A VGND VGND VPWR VPWR _14035_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ _13298_/CLK _12687_/D VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__dfxtp_1
X_14426_ _14732_/CLK _14426_/D VGND VGND VPWR VPWR _14426_/Q sky130_fd_sc_hd__dfxtp_1
X_11638_ _11638_/A VGND VGND VPWR VPWR _13994_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14357_ _14357_/CLK _14357_/D VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__dfxtp_1
XFILLER_144_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11569_ _11569_/A VGND VGND VPWR VPWR _13866_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13308_ _13570_/CLK hold413/X VGND VGND VPWR VPWR _13308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14288_ _14292_/CLK _14288_/D VGND VGND VPWR VPWR _14288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13239_ _14010_/CLK _13746_/Q VGND VGND VPWR VPWR _13511_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_112_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07800_ _07797_/Y _13169_/D _07800_/S VGND VGND VPWR VPWR _07801_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08780_ _13464_/Q _09569_/B VGND VGND VPWR VPWR _08780_/X sky130_fd_sc_hd__or2_1
XFILLER_97_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05992_ _05992_/A _05992_/B _05992_/C VGND VGND VPWR VPWR _05993_/D sky130_fd_sc_hd__and3_1
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07731_ _07731_/A _07757_/B VGND VGND VPWR VPWR _07732_/B sky130_fd_sc_hd__xnor2_1
XFILLER_78_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07662_ _07637_/Y _07661_/Y _11266_/A VGND VGND VPWR VPWR _07663_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06613_ _06613_/A _06613_/B VGND VGND VPWR VPWR _12903_/D sky130_fd_sc_hd__nor2_1
X_09401_ _13594_/Q _09401_/B VGND VGND VPWR VPWR _09401_/Y sky130_fd_sc_hd__nor2_1
X_07593_ _07645_/A VGND VGND VPWR VPWR _07622_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09332_ _13303_/Q _13541_/Q _09332_/S VGND VGND VPWR VPWR _09333_/A sky130_fd_sc_hd__mux2_1
X_06544_ _10337_/B _06544_/B _06563_/B VGND VGND VPWR VPWR _06552_/B sky130_fd_sc_hd__and3_1
XFILLER_33_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09263_ _13550_/Q _09270_/B VGND VGND VPWR VPWR _09267_/B sky130_fd_sc_hd__xnor2_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06475_ _06449_/A _06463_/A _06462_/X VGND VGND VPWR VPWR _06475_/Y sky130_fd_sc_hd__o21ai_1
X_08214_ _08223_/A _08214_/B VGND VGND VPWR VPWR _08214_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_21_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09194_ _13539_/Q _09206_/B VGND VGND VPWR VPWR _09220_/A sky130_fd_sc_hd__xnor2_1
XFILLER_21_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08145_ _08228_/S _08141_/X _08144_/X _08208_/A VGND VGND VPWR VPWR _08145_/X sky130_fd_sc_hd__o211a_1
XFILLER_147_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08076_ _12974_/Q _13274_/Q _08084_/S VGND VGND VPWR VPWR _08077_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07027_ _07040_/A _07139_/A _07045_/C VGND VGND VPWR VPWR _07028_/B sky130_fd_sc_hd__a21oi_1
XFILLER_161_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08978_ _08978_/A _08978_/B _08991_/C _08978_/D VGND VGND VPWR VPWR _08979_/B sky130_fd_sc_hd__and4_1
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_152_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_152_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold67 hold67/A VGND VGND VPWR VPWR hold67/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold78 hold78/A VGND VGND VPWR VPWR hold78/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_07929_ _13269_/Q _07962_/B VGND VGND VPWR VPWR _07930_/B sky130_fd_sc_hd__or2_1
XFILLER_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold89 hold89/A VGND VGND VPWR VPWR hold89/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_10940_ _12586_/A VGND VGND VPWR VPWR _10940_/X sky130_fd_sc_hd__buf_2
XFILLER_56_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10871_ _10871_/A VGND VGND VPWR VPWR _13194_/D sky130_fd_sc_hd__clkbuf_1
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12610_ _14733_/Q _12608_/B _12609_/X VGND VGND VPWR VPWR _12611_/B sky130_fd_sc_hd__o21ai_1
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13590_ _14012_/CLK _13590_/D repeater56/X VGND VGND VPWR VPWR _13590_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12541_ _11323_/X _14716_/Q _12543_/S VGND VGND VPWR VPWR _12542_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12472_ _14667_/Q _12013_/A _12472_/S VGND VGND VPWR VPWR _12473_/A sky130_fd_sc_hd__mux2_1
X_14211_ _14212_/CLK _14211_/D VGND VGND VPWR VPWR _14211_/Q sky130_fd_sc_hd__dfxtp_1
X_11423_ _13734_/Q _11427_/B VGND VGND VPWR VPWR _11424_/A sky130_fd_sc_hd__and2_1
XFILLER_126_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 hold42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11354_ _12013_/A VGND VGND VPWR VPWR _11354_/X sky130_fd_sc_hd__clkbuf_2
X_14142_ _14294_/CLK _14142_/D VGND VGND VPWR VPWR _14142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10305_ _10306_/A _13511_/D _10306_/C VGND VGND VPWR VPWR _10307_/A sky130_fd_sc_hd__o21a_1
X_11285_ _14695_/Q VGND VGND VPWR VPWR _11285_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14073_ _14726_/CLK _14073_/D VGND VGND VPWR VPWR _14073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10236_ _14521_/D _10236_/B VGND VGND VPWR VPWR _10237_/B sky130_fd_sc_hd__nor2_1
X_13024_ _13027_/CLK _13024_/D repeater59/X VGND VGND VPWR VPWR _13024_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10167_ _10167_/A VGND VGND VPWR VPWR _14134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10098_ _10139_/A _14142_/Q VGND VGND VPWR VPWR _10182_/S sky130_fd_sc_hd__xor2_2
X_13926_ _14196_/CLK hold93/X VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13857_ _14179_/CLK _13857_/D VGND VGND VPWR VPWR _13857_/Q sky130_fd_sc_hd__dfxtp_1
X_12808_ _13622_/CLK _12808_/D VGND VGND VPWR VPWR hold329/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13788_ _13799_/CLK _13788_/D VGND VGND VPWR VPWR _13788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12739_ _14333_/CLK _12739_/D VGND VGND VPWR VPWR hold420/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06260_ _13955_/Q _13947_/Q _10023_/A VGND VGND VPWR VPWR _06260_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14409_ _14425_/CLK _14409_/D VGND VGND VPWR VPWR hold281/A sky130_fd_sc_hd__dfxtp_1
X_06191_ _06191_/A VGND VGND VPWR VPWR _14365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold504 hold504/A VGND VGND VPWR VPWR hold504/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold515 hold515/A VGND VGND VPWR VPWR hold515/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09950_ _09950_/A VGND VGND VPWR VPWR _12861_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08901_ _08901_/A _08901_/B VGND VGND VPWR VPWR _08903_/A sky130_fd_sc_hd__xnor2_1
XFILLER_103_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _13691_/Q _13692_/Q _13693_/Q _09881_/D VGND VGND VPWR VPWR _09885_/B sky130_fd_sc_hd__and4_1
XFILLER_97_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08832_ _08851_/B _08907_/B _08929_/A _08907_/A VGND VGND VPWR VPWR _08832_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_111_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05975_ _13629_/Q _13638_/Q _13639_/Q _13640_/Q VGND VGND VPWR VPWR _05976_/C sky130_fd_sc_hd__or4_1
X_08763_ _08770_/A _08763_/B _08763_/C VGND VGND VPWR VPWR _08763_/Y sky130_fd_sc_hd__nand3_1
X_07714_ _07683_/A _07683_/B _07713_/Y VGND VGND VPWR VPWR _07715_/B sky130_fd_sc_hd__o21bai_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ _08698_/A _08714_/B VGND VGND VPWR VPWR _08694_/X sky130_fd_sc_hd__or2_1
XFILLER_53_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07645_ _07645_/A _07645_/B _13246_/D _07723_/C VGND VGND VPWR VPWR _07688_/A sky130_fd_sc_hd__and4_1
XFILLER_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07576_ _07570_/X _07573_/Y _07574_/X _07575_/X VGND VGND VPWR VPWR _13160_/D sky130_fd_sc_hd__a31o_1
XFILLER_22_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09315_ _13295_/Q _13533_/Q _09321_/S VGND VGND VPWR VPWR _09316_/A sky130_fd_sc_hd__mux2_1
X_06527_ _06527_/A VGND VGND VPWR VPWR _06527_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06458_ _14436_/Q _14434_/Q _06458_/S VGND VGND VPWR VPWR _06458_/X sky130_fd_sc_hd__mux2_1
X_09246_ _13547_/Q _09250_/B VGND VGND VPWR VPWR _09255_/A sky130_fd_sc_hd__xor2_1
X_09177_ _09177_/A _09177_/B VGND VGND VPWR VPWR _09177_/X sky130_fd_sc_hd__or2_1
X_06389_ _12910_/Q VGND VGND VPWR VPWR _06622_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08128_ _08142_/A _14003_/Q VGND VGND VPWR VPWR _08128_/X sky130_fd_sc_hd__and2b_1
XFILLER_107_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08059_ _08059_/A VGND VGND VPWR VPWR _12690_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput35 _13332_/Q VGND VGND VPWR VPWR data_o[14] sky130_fd_sc_hd__buf_2
XFILLER_122_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput46 _13320_/Q VGND VGND VPWR VPWR data_o[2] sky130_fd_sc_hd__buf_2
XFILLER_89_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11070_ _11070_/A _11013_/X VGND VGND VPWR VPWR _11070_/X sky130_fd_sc_hd__or2b_1
XFILLER_1_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10021_ _13911_/D _13978_/Q _13910_/D _06047_/X _13976_/Q VGND VGND VPWR VPWR _13924_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11972_ _14700_/Q VGND VGND VPWR VPWR _11972_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13711_ _14251_/CLK _13711_/D VGND VGND VPWR VPWR _13711_/Q sky130_fd_sc_hd__dfxtp_1
X_10923_ _14013_/Q _13979_/Q _13819_/Q _14531_/Q _10921_/X _10922_/X VGND VGND VPWR
+ VPWR _10926_/A sky130_fd_sc_hd__mux4_1
XFILLER_44_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14691_ _14710_/CLK hold82/X VGND VGND VPWR VPWR hold309/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13642_ _13653_/CLK hold325/X VGND VGND VPWR VPWR _13642_/Q sky130_fd_sc_hd__dfxtp_1
X_10854_ _10876_/A VGND VGND VPWR VPWR _10863_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_32_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13573_ _14098_/CLK hold167/X VGND VGND VPWR VPWR _13573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10785_ _10785_/A VGND VGND VPWR VPWR _13055_/D sky130_fd_sc_hd__clkbuf_1
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12524_ _11297_/X _14708_/Q _12532_/S VGND VGND VPWR VPWR _12525_/A sky130_fd_sc_hd__mux2_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12455_ _14659_/Q _14516_/Q _12461_/S VGND VGND VPWR VPWR _12456_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11406_ _11406_/A VGND VGND VPWR VPWR _13795_/D sky130_fd_sc_hd__clkbuf_1
X_12386_ _14615_/Q _12013_/X _12386_/S VGND VGND VPWR VPWR _12387_/A sky130_fd_sc_hd__mux2_1
X_14125_ _14608_/CLK hold56/X VGND VGND VPWR VPWR _14125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11337_ _12004_/A VGND VGND VPWR VPWR _11337_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14056_ _14539_/CLK _14056_/D VGND VGND VPWR VPWR _14056_/Q sky130_fd_sc_hd__dfxtp_1
X_11268_ _11268_/A _11268_/B VGND VGND VPWR VPWR _11269_/A sky130_fd_sc_hd__and2_1
X_13007_ _13296_/CLK _13007_/D hold1/X VGND VGND VPWR VPWR _13007_/Q sky130_fd_sc_hd__dfrtp_1
X_10219_ _10219_/A VGND VGND VPWR VPWR _14397_/D sky130_fd_sc_hd__clkbuf_1
X_11199_ _11136_/X _11196_/X _11198_/X _11157_/X VGND VGND VPWR VPWR _11199_/X sky130_fd_sc_hd__o211a_1
XFILLER_94_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13909_ _14179_/CLK _13909_/D VGND VGND VPWR VPWR _13909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07430_ _13144_/Q _07435_/A _07435_/B VGND VGND VPWR VPWR _07438_/A sky130_fd_sc_hd__and3_1
XFILLER_51_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07361_ _07387_/A _07361_/B VGND VGND VPWR VPWR _07374_/A sky130_fd_sc_hd__or2_1
XFILLER_149_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06312_ _06312_/A VGND VGND VPWR VPWR _14190_/D sky130_fd_sc_hd__clkbuf_1
X_09100_ _09109_/A _09099_/X VGND VGND VPWR VPWR _09103_/A sky130_fd_sc_hd__or2b_1
X_07292_ _13133_/Q _09101_/B VGND VGND VPWR VPWR _07292_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09031_ _09655_/S VGND VGND VPWR VPWR _09040_/S sky130_fd_sc_hd__clkbuf_2
X_06243_ _14092_/Q _06245_/B VGND VGND VPWR VPWR _06244_/A sky130_fd_sc_hd__and2_1
XFILLER_164_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06174_ _06174_/A VGND VGND VPWR VPWR _14174_/D sky130_fd_sc_hd__clkbuf_1
Xhold301 hold301/A VGND VGND VPWR VPWR hold301/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold312 hold312/A VGND VGND VPWR VPWR hold312/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold323 hold323/A VGND VGND VPWR VPWR hold323/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold334 hold334/A VGND VGND VPWR VPWR hold334/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14752__63 VGND VGND VPWR VPWR _14752__63/HI data_o[26] sky130_fd_sc_hd__conb_1
Xhold345 hold345/A VGND VGND VPWR VPWR hold345/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold356 hold356/A VGND VGND VPWR VPWR hold356/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold367 hold367/A VGND VGND VPWR VPWR hold367/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_117_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold378 hold378/A VGND VGND VPWR VPWR hold378/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold389 hold389/A VGND VGND VPWR VPWR hold389/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09933_ _13491_/Q _13680_/Q _09935_/S VGND VGND VPWR VPWR _09934_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _13687_/Q _09870_/B _09776_/X VGND VGND VPWR VPWR _09865_/B sky130_fd_sc_hd__o21ai_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ _08828_/A _08927_/A _08833_/C VGND VGND VPWR VPWR _08816_/B sky130_fd_sc_hd__a21oi_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09795_ _09795_/A _09795_/B VGND VGND VPWR VPWR _09796_/B sky130_fd_sc_hd__and2_1
X_08746_ _08746_/A VGND VGND VPWR VPWR _09542_/B sky130_fd_sc_hd__buf_2
X_05958_ _13635_/Q _13636_/Q _13637_/Q _13642_/Q VGND VGND VPWR VPWR _05959_/D sky130_fd_sc_hd__and4_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _09525_/B VGND VGND VPWR VPWR _08746_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ _07613_/A _07745_/A _07626_/Y _07656_/A VGND VGND VPWR VPWR _07641_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07559_ _07559_/A _07559_/B VGND VGND VPWR VPWR _07559_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10570_ _10570_/A _10570_/B _10570_/C VGND VGND VPWR VPWR _10571_/B sky130_fd_sc_hd__nand3_1
XFILLER_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09229_ _09229_/A _09228_/X VGND VGND VPWR VPWR _09242_/C sky130_fd_sc_hd__or2b_1
X_12240_ _11297_/X _14536_/Q _12248_/S VGND VGND VPWR VPWR _12241_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12171_ _12171_/A VGND VGND VPWR VPWR _14497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11122_ _11088_/X _11118_/Y _11121_/Y _11095_/X VGND VGND VPWR VPWR _11123_/B sky130_fd_sc_hd__a211o_1
XFILLER_111_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11053_ _13325_/Q _11008_/X _11042_/X _11052_/Y VGND VGND VPWR VPWR _13325_/D sky130_fd_sc_hd__o22a_1
XFILLER_77_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10004_ _14628_/Q _14626_/Q _14647_/Q VGND VGND VPWR VPWR _10004_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14743_ _14749_/CLK _14743_/D VGND VGND VPWR VPWR _14743_/Q sky130_fd_sc_hd__dfxtp_1
X_11955_ _11955_/A VGND VGND VPWR VPWR _14295_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10906_ _11185_/A VGND VGND VPWR VPWR _12626_/B sky130_fd_sc_hd__buf_2
X_14674_ _14687_/CLK _14674_/D VGND VGND VPWR VPWR hold267/A sky130_fd_sc_hd__dfxtp_1
XFILLER_60_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11886_ _14240_/Q _11510_/X _11886_/S VGND VGND VPWR VPWR _11887_/A sky130_fd_sc_hd__mux2_1
X_13625_ _13635_/CLK hold385/X VGND VGND VPWR VPWR _13625_/Q sky130_fd_sc_hd__dfxtp_1
X_10837_ _13137_/Q _10841_/B VGND VGND VPWR VPWR _10838_/A sky130_fd_sc_hd__and2_1
XFILLER_13_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13556_ _13558_/CLK hold163/X VGND VGND VPWR VPWR _13556_/Q sky130_fd_sc_hd__dfxtp_1
X_10768_ _13006_/Q _10768_/B VGND VGND VPWR VPWR _10769_/A sky130_fd_sc_hd__and2_1
X_12507_ _12506_/Y _14157_/Q _14110_/Q VGND VGND VPWR VPWR _14693_/D sky130_fd_sc_hd__a21o_1
XFILLER_157_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13487_ _13721_/CLK hold176/X VGND VGND VPWR VPWR _13487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10699_ _10699_/A VGND VGND VPWR VPWR _12928_/D sky130_fd_sc_hd__clkbuf_1
X_12438_ _12438_/A VGND VGND VPWR VPWR _14651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12369_ _14607_/Q _11988_/X _12375_/S VGND VGND VPWR VPWR _12370_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14108_ _14108_/CLK _14108_/D VGND VGND VPWR VPWR _14108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14039_ _14047_/CLK _14039_/D VGND VGND VPWR VPWR _14039_/Q sky130_fd_sc_hd__dfxtp_1
X_06930_ _07940_/A VGND VGND VPWR VPWR _06930_/X sky130_fd_sc_hd__buf_2
XFILLER_110_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06861_ _07802_/A VGND VGND VPWR VPWR _06861_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08600_ _08590_/B _08621_/B _08621_/A VGND VGND VPWR VPWR _08601_/B sky130_fd_sc_hd__a21o_1
X_09580_ _09502_/X _09578_/X _09579_/Y _09506_/X VGND VGND VPWR VPWR _13619_/D sky130_fd_sc_hd__a31o_1
X_06792_ _06794_/A _06794_/B _06827_/B VGND VGND VPWR VPWR _06793_/B sky130_fd_sc_hd__a21o_1
XFILLER_36_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08531_ _08531_/A _08531_/B VGND VGND VPWR VPWR _08531_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_51_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08462_ _08462_/A VGND VGND VPWR VPWR _13436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07413_ _07414_/C _07412_/X VGND VGND VPWR VPWR _07425_/B sky130_fd_sc_hd__or2b_1
XFILLER_50_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08393_ _13093_/Q _13374_/Q _08395_/S VGND VGND VPWR VPWR _08394_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07344_ _13169_/Q _13666_/Q _07344_/S VGND VGND VPWR VPWR _07344_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07275_ _13133_/Q _09101_/B VGND VGND VPWR VPWR _07276_/C sky130_fd_sc_hd__and2_1
XFILLER_149_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06226_ _14400_/Q _14392_/Q _06321_/S VGND VGND VPWR VPWR _06226_/X sky130_fd_sc_hd__mux2_1
X_09014_ _13208_/Q _13437_/Q _09018_/S VGND VGND VPWR VPWR _09015_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06157_ _10616_/B _06156_/X _10121_/S VGND VGND VPWR VPWR _06158_/A sky130_fd_sc_hd__mux2_1
Xhold120 hold120/A VGND VGND VPWR VPWR hold120/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold131 hold131/A VGND VGND VPWR VPWR hold131/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold142 hold142/A VGND VGND VPWR VPWR hold142/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold153 hold153/A VGND VGND VPWR VPWR hold153/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold164 hold164/A VGND VGND VPWR VPWR hold164/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06088_ _06088_/A VGND VGND VPWR VPWR _13967_/D sky130_fd_sc_hd__clkbuf_1
Xhold175 hold175/A VGND VGND VPWR VPWR hold175/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold186 hold186/A VGND VGND VPWR VPWR hold186/X sky130_fd_sc_hd__clkbuf_2
Xhold197 hold197/A VGND VGND VPWR VPWR hold197/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09916_ _13483_/Q _13672_/Q _09924_/S VGND VGND VPWR VPWR _09917_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09847_ _09858_/C VGND VGND VPWR VPWR _09851_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _09778_/A _09778_/B _09778_/C VGND VGND VPWR VPWR _09785_/B sky130_fd_sc_hd__and3_1
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _13457_/Q _09525_/B VGND VGND VPWR VPWR _08739_/A sky130_fd_sc_hd__and2_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11740_/A VGND VGND VPWR VPWR _14061_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _11671_/A VGND VGND VPWR VPWR _14018_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13410_ _13617_/CLK hold468/X VGND VGND VPWR VPWR _13410_/Q sky130_fd_sc_hd__dfxtp_1
X_10622_ _14294_/Q _10620_/X _10621_/X _14293_/Q _14282_/Q VGND VGND VPWR VPWR _14289_/D
+ sky130_fd_sc_hd__a221o_1
X_14390_ _14410_/CLK _14390_/D VGND VGND VPWR VPWR _14390_/Q sky130_fd_sc_hd__dfxtp_1
X_13341_ _14619_/CLK _13341_/D VGND VGND VPWR VPWR _13341_/Q sky130_fd_sc_hd__dfxtp_1
X_10553_ _10553_/A _10553_/B VGND VGND VPWR VPWR _10562_/B sky130_fd_sc_hd__nor2_1
XFILLER_154_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13272_ _13273_/CLK _13272_/D repeater59/X VGND VGND VPWR VPWR _13272_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10484_ _10444_/B _10501_/C _10485_/C VGND VGND VPWR VPWR _10486_/A sky130_fd_sc_hd__a21oi_1
X_12223_ _12223_/A VGND VGND VPWR VPWR _14518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12154_ _12154_/A VGND VGND VPWR VPWR _14489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11105_ _14268_/Q _14659_/Q _13766_/Q _14714_/Q _11091_/X _11092_/X VGND VGND VPWR
+ VPWR _11106_/B sky130_fd_sc_hd__mux4_1
XFILLER_78_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12085_ _11354_/X _14460_/Q _12085_/S VGND VGND VPWR VPWR _12086_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11036_ _11017_/X _11033_/Y _11035_/Y _11024_/X VGND VGND VPWR VPWR _11037_/B sky130_fd_sc_hd__a211o_1
XFILLER_64_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12987_ _14636_/CLK _12987_/D VGND VGND VPWR VPWR _13108_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_80_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14726_ _14726_/CLK _14726_/D VGND VGND VPWR VPWR _14726_/Q sky130_fd_sc_hd__dfxtp_1
X_11938_ _14275_/Q _11507_/X _11940_/S VGND VGND VPWR VPWR _11939_/A sky130_fd_sc_hd__mux2_1
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14657_ _14657_/CLK _14657_/D VGND VGND VPWR VPWR _14657_/Q sky130_fd_sc_hd__dfxtp_1
X_11869_ _14232_/Q _11485_/X _11875_/S VGND VGND VPWR VPWR _11870_/A sky130_fd_sc_hd__mux2_1
X_13608_ _13610_/CLK _13608_/D repeater57/X VGND VGND VPWR VPWR _13608_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_159_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14588_ _14588_/CLK hold101/X VGND VGND VPWR VPWR _14588_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13539_ _13558_/CLK _13539_/D _12609_/A VGND VGND VPWR VPWR _13539_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_146_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07060_ _13708_/Q VGND VGND VPWR VPWR _07141_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06011_ _13563_/Q _13572_/Q _13573_/Q _13574_/Q VGND VGND VPWR VPWR _06012_/C sky130_fd_sc_hd__and4_1
XFILLER_126_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07962_ _13274_/Q _07962_/B VGND VGND VPWR VPWR _07970_/A sky130_fd_sc_hd__and2_1
XFILLER_102_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09701_ _09715_/S _14440_/Q _09718_/A VGND VGND VPWR VPWR _09701_/X sky130_fd_sc_hd__a21o_1
X_06913_ _06914_/A _06914_/B _06924_/C VGND VGND VPWR VPWR _06919_/B sky130_fd_sc_hd__a21o_1
X_07893_ _07893_/A _07893_/B _07893_/C VGND VGND VPWR VPWR _07893_/Y sky130_fd_sc_hd__nand3_1
XFILLER_28_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09632_ _09632_/A VGND VGND VPWR VPWR _12829_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06844_ _13011_/Q _07895_/B _07895_/C VGND VGND VPWR VPWR _06851_/A sky130_fd_sc_hd__and3_1
XFILLER_28_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09563_ _13617_/Q _09563_/B VGND VGND VPWR VPWR _09564_/B sky130_fd_sc_hd__nor2_1
X_06775_ _06775_/A _06775_/B VGND VGND VPWR VPWR _06775_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08514_ _08733_/A VGND VGND VPWR VPWR _08665_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09494_ _08504_/X _09492_/X _09493_/X VGND VGND VPWR VPWR _13606_/D sky130_fd_sc_hd__a21o_1
XFILLER_24_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08445_ _14248_/Q _14246_/Q _08472_/A VGND VGND VPWR VPWR _08445_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08376_ _13085_/Q _13366_/Q _08384_/S VGND VGND VPWR VPWR _08377_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07327_ _07327_/A VGND VGND VPWR VPWR _07327_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07258_ _07258_/A _07258_/B VGND VGND VPWR VPWR _07258_/Y sky130_fd_sc_hd__nand2_1
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06209_ _14408_/Q _14400_/Q hold94/A VGND VGND VPWR VPWR _06324_/A sky130_fd_sc_hd__mux2_1
X_07189_ _07190_/B _07203_/C _07203_/B _07190_/A VGND VGND VPWR VPWR _07191_/A sky130_fd_sc_hd__a22oi_1
XFILLER_105_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12910_ _13263_/CLK hold505/X VGND VGND VPWR VPWR _12910_/Q sky130_fd_sc_hd__dfxtp_2
X_13890_ _14657_/CLK hold371/X VGND VGND VPWR VPWR _13890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12841_ _13721_/CLK _12841_/D VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12772_ _13698_/CLK _12772_/D VGND VGND VPWR VPWR hold263/A sky130_fd_sc_hd__dfxtp_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14619_/CLK _14511_/D VGND VGND VPWR VPWR _14511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11291_/X _14054_/Q _11725_/S VGND VGND VPWR VPWR _11724_/A sky130_fd_sc_hd__mux2_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14442_ _14704_/CLK _14442_/D VGND VGND VPWR VPWR _14442_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _11654_/A VGND VGND VPWR VPWR _14002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10605_ _10603_/X _10604_/X _13886_/Q VGND VGND VPWR VPWR _13885_/D sky130_fd_sc_hd__o21a_1
X_14373_ _14536_/CLK _14373_/D VGND VGND VPWR VPWR hold366/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11585_ _13650_/Q _11585_/B VGND VGND VPWR VPWR _11586_/A sky130_fd_sc_hd__and2_1
XFILLER_155_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13324_ _14709_/CLK _13324_/D VGND VGND VPWR VPWR _13324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10536_ _10549_/A _10536_/B VGND VGND VPWR VPWR _10537_/B sky130_fd_sc_hd__nand2_1
XFILLER_128_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13255_ _13258_/CLK _13255_/D hold1/X VGND VGND VPWR VPWR _13255_/Q sky130_fd_sc_hd__dfrtp_1
X_10467_ _10468_/A _10468_/B VGND VGND VPWR VPWR _10469_/A sky130_fd_sc_hd__and2_1
XFILLER_142_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12206_ _14120_/Q _14117_/Q _12205_/X VGND VGND VPWR VPWR _12206_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_142_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13186_ _13423_/CLK _13186_/D VGND VGND VPWR VPWR hold358/A sky130_fd_sc_hd__dfxtp_1
XFILLER_124_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10398_ _10378_/X _10398_/B VGND VGND VPWR VPWR _10411_/B sky130_fd_sc_hd__and2b_1
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12137_ _14483_/Q _12010_/X _12139_/S VGND VGND VPWR VPWR _12138_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12068_ _11317_/X _14452_/Q _12074_/S VGND VGND VPWR VPWR _12069_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11019_ _11019_/A VGND VGND VPWR VPWR _11019_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06560_ _06567_/A _06560_/B VGND VGND VPWR VPWR _06560_/Y sky130_fd_sc_hd__xnor2_1
X_14709_ _14709_/CLK _14709_/D VGND VGND VPWR VPWR _14709_/Q sky130_fd_sc_hd__dfxtp_1
X_06491_ _06486_/B _06490_/Y _06530_/S VGND VGND VPWR VPWR _06492_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08230_ _08250_/C VGND VGND VPWR VPWR _08279_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08161_ _14008_/Q _14006_/Q _08161_/S VGND VGND VPWR VPWR _08161_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07112_ _13707_/Q hold177/A VGND VGND VPWR VPWR _07113_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08092_ _08092_/A VGND VGND VPWR VPWR _12705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07043_ _13706_/Q VGND VGND VPWR VPWR _07119_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08994_ _08994_/A _08994_/B VGND VGND VPWR VPWR _08995_/B sky130_fd_sc_hd__nor2_1
XFILLER_142_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07945_ _07909_/X _07943_/X _07944_/Y _07940_/X VGND VGND VPWR VPWR _13271_/D sky130_fd_sc_hd__a31o_1
XFILLER_68_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07876_ _13262_/Q _07876_/B VGND VGND VPWR VPWR _07881_/A sky130_fd_sc_hd__nand2_1
X_09615_ _09615_/A VGND VGND VPWR VPWR _12821_/D sky130_fd_sc_hd__clkbuf_1
X_06827_ _06827_/A _06827_/B VGND VGND VPWR VPWR _06827_/X sky130_fd_sc_hd__or2_1
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09546_ _13613_/Q _13614_/Q _08787_/B VGND VGND VPWR VPWR _09553_/B sky130_fd_sc_hd__o21ai_1
X_06758_ _13005_/Q _07846_/B _07846_/C VGND VGND VPWR VPWR _06775_/B sky130_fd_sc_hd__and3_1
XFILLER_70_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09477_ _09477_/A _09477_/B VGND VGND VPWR VPWR _09478_/B sky130_fd_sc_hd__nor2_1
X_06689_ _06636_/Y _06812_/B _06688_/X _06634_/X VGND VGND VPWR VPWR _06689_/X sky130_fd_sc_hd__a22o_1
X_08428_ _13475_/Q VGND VGND VPWR VPWR _08470_/A sky130_fd_sc_hd__inv_2
XFILLER_7_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08359_ _08359_/A VGND VGND VPWR VPWR _12713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11370_ _12022_/A VGND VGND VPWR VPWR _11370_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_137_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10321_ _13746_/Q _13106_/Q _10321_/C VGND VGND VPWR VPWR _10322_/B sky130_fd_sc_hd__nor3_1
XFILLER_164_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13040_ _14636_/CLK _13040_/D VGND VGND VPWR VPWR hold180/A sky130_fd_sc_hd__dfxtp_1
X_10252_ _10238_/X _10251_/X _14556_/D VGND VGND VPWR VPWR _10252_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10183_ _10183_/A VGND VGND VPWR VPWR _14139_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13942_ _13972_/CLK _13942_/D VGND VGND VPWR VPWR _13942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13873_ _14656_/CLK _13873_/D VGND VGND VPWR VPWR _13873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12824_ _13653_/CLK _12824_/D VGND VGND VPWR VPWR hold337/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ _13704_/CLK _12755_/D VGND VGND VPWR VPWR hold169/A sky130_fd_sc_hd__dfxtp_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _14035_/Q _11519_/X _11708_/S VGND VGND VPWR VPWR _11707_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _13298_/CLK _12686_/D VGND VGND VPWR VPWR hold240/A sky130_fd_sc_hd__dfxtp_1
X_14425_ _14425_/CLK _14425_/D VGND VGND VPWR VPWR _14425_/Q sky130_fd_sc_hd__dfxtp_1
X_11637_ _13994_/Q _11497_/X _11645_/S VGND VGND VPWR VPWR _11638_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14356_ _14357_/CLK _14356_/D VGND VGND VPWR VPWR hold472/A sky130_fd_sc_hd__dfxtp_1
X_11568_ _13642_/Q _11574_/B VGND VGND VPWR VPWR _11569_/A sky130_fd_sc_hd__and2_1
XFILLER_116_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13307_ _13570_/CLK hold193/X VGND VGND VPWR VPWR _13307_/Q sky130_fd_sc_hd__dfxtp_1
X_10519_ _10519_/A _10526_/C VGND VGND VPWR VPWR _10539_/A sky130_fd_sc_hd__and2_1
XFILLER_6_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14287_ _14292_/CLK _14287_/D VGND VGND VPWR VPWR _14287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11499_ _13834_/Q _11497_/X _11511_/S VGND VGND VPWR VPWR _11500_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13238_ _13621_/CLK hold80/X VGND VGND VPWR VPWR _13238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13169_ _13666_/CLK _13169_/D VGND VGND VPWR VPWR _13169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05991_ _14099_/Q _14100_/Q _14101_/Q _14102_/Q VGND VGND VPWR VPWR _05992_/C sky130_fd_sc_hd__and4_1
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07730_ _07697_/A _07697_/B _07703_/A _07703_/B VGND VGND VPWR VPWR _07757_/B sky130_fd_sc_hd__a22o_1
XFILLER_111_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07661_ _07738_/A _07661_/B VGND VGND VPWR VPWR _07661_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_1_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09400_ _13594_/Q _09401_/B VGND VGND VPWR VPWR _09400_/Y sky130_fd_sc_hd__nand2_1
X_06612_ _12903_/Q _06620_/B _06599_/X VGND VGND VPWR VPWR _06613_/B sky130_fd_sc_hd__o21ai_1
X_07592_ _13110_/Q VGND VGND VPWR VPWR _07645_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09331_ _09331_/A VGND VGND VPWR VPWR _12792_/D sky130_fd_sc_hd__clkbuf_1
X_06543_ _06543_/A VGND VGND VPWR VPWR _10337_/B sky130_fd_sc_hd__buf_2
XFILLER_33_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09262_ _08218_/X _09264_/B _09261_/Y _09215_/X VGND VGND VPWR VPWR _13549_/D sky130_fd_sc_hd__a31o_1
X_06474_ _06493_/A _06474_/B VGND VGND VPWR VPWR _06488_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08213_ _08193_/A _08193_/B _08204_/A _08212_/Y VGND VGND VPWR VPWR _08214_/B sky130_fd_sc_hd__o31ai_2
X_09193_ _09186_/A _09188_/Y _09190_/Y _09173_/B _09192_/Y VGND VGND VPWR VPWR _09195_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_119_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08144_ _08197_/A _13477_/Q _08176_/A VGND VGND VPWR VPWR _08144_/X sky130_fd_sc_hd__a21o_1
XFILLER_146_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08075_ _08097_/A VGND VGND VPWR VPWR _08084_/S sky130_fd_sc_hd__buf_2
XFILLER_161_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07026_ _07063_/A _07139_/A _07045_/C VGND VGND VPWR VPWR _07028_/A sky130_fd_sc_hd__and3_1
XFILLER_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_08977_ _08978_/B _08991_/C _08991_/B _08978_/A VGND VGND VPWR VPWR _08979_/A sky130_fd_sc_hd__a22oi_1
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_07928_ _13269_/Q _07963_/B VGND VGND VPWR VPWR _07939_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold68 hold68/A VGND VGND VPWR VPWR hold68/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold79 hold79/A VGND VGND VPWR VPWR hold79/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07859_ _07859_/A _07859_/B _07859_/C _07859_/D VGND VGND VPWR VPWR _07860_/B sky130_fd_sc_hd__nor4_2
XFILLER_71_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10870_ _13152_/Q _10874_/B VGND VGND VPWR VPWR _10871_/A sky130_fd_sc_hd__and2_1
XFILLER_72_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09529_ _09532_/B _09528_/X _08735_/X VGND VGND VPWR VPWR _13611_/D sky130_fd_sc_hd__o21bai_1
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12540_ _12540_/A VGND VGND VPWR VPWR _14715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12471_ _12471_/A VGND VGND VPWR VPWR _14666_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14210_ _14210_/CLK _14210_/D VGND VGND VPWR VPWR _14210_/Q sky130_fd_sc_hd__dfxtp_1
X_11422_ _11422_/A VGND VGND VPWR VPWR _13802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14141_ _14159_/CLK _14141_/D VGND VGND VPWR VPWR _14141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11353_ _11362_/C _11353_/B _11353_/C VGND VGND VPWR VPWR _12013_/A sky130_fd_sc_hd__and3b_4
XFILLER_152_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10304_ _10304_/A _13512_/D VGND VGND VPWR VPWR _10306_/C sky130_fd_sc_hd__xor2_1
XFILLER_141_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14072_ _14617_/CLK _14072_/D VGND VGND VPWR VPWR _14072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11284_ _11284_/A VGND VGND VPWR VPWR _13755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13023_ _13027_/CLK _13023_/D repeater59/X VGND VGND VPWR VPWR _13023_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_140_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10235_ _14367_/Q _10230_/X _10237_/A VGND VGND VPWR VPWR _14524_/D sky130_fd_sc_hd__a21o_1
XFILLER_79_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10166_ _10161_/X _10165_/X _14292_/D VGND VGND VPWR VPWR _10167_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10097_ _14141_/Q VGND VGND VPWR VPWR _10139_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_35_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13925_ _14050_/CLK hold39/X VGND VGND VPWR VPWR _13925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13856_ _14180_/CLK _13856_/D VGND VGND VPWR VPWR _13856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12807_ _14530_/CLK _12807_/D VGND VGND VPWR VPWR hold476/A sky130_fd_sc_hd__dfxtp_1
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13787_ _13799_/CLK _13787_/D VGND VGND VPWR VPWR _13787_/Q sky130_fd_sc_hd__dfxtp_1
X_10999_ _10991_/X _10996_/X _10998_/X _10929_/X VGND VGND VPWR VPWR _10999_/X sky130_fd_sc_hd__o211a_1
XFILLER_43_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _14333_/CLK _12738_/D VGND VGND VPWR VPWR hold98/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12669_ _13351_/CLK _12669_/D VGND VGND VPWR VPWR _12991_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_129_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14408_ _14410_/CLK _14408_/D VGND VGND VPWR VPWR _14408_/Q sky130_fd_sc_hd__dfxtp_1
X_06190_ _06186_/X _06187_/X _06197_/A VGND VGND VPWR VPWR _06191_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14339_ _14697_/CLK hold478/X VGND VGND VPWR VPWR _14339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold505 hold505/A VGND VGND VPWR VPWR hold505/X sky130_fd_sc_hd__clkbuf_1
Xhold516 hold516/A VGND VGND VPWR VPWR hold516/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08900_ _13518_/D _13430_/Q VGND VGND VPWR VPWR _08901_/B sky130_fd_sc_hd__nand2_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _13692_/Q _09878_/A _09879_/Y VGND VGND VPWR VPWR _13692_/D sky130_fd_sc_hd__a21oi_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _13517_/D VGND VGND VPWR VPWR _08907_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _08763_/B _08763_/C _08770_/A VGND VGND VPWR VPWR _08767_/B sky130_fd_sc_hd__a21o_1
X_05974_ _13641_/Q _13646_/Q _13647_/Q _13648_/Q VGND VGND VPWR VPWR _05976_/B sky130_fd_sc_hd__or4_1
XFILLER_66_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07713_ _07713_/A _07713_/B VGND VGND VPWR VPWR _07713_/Y sky130_fd_sc_hd__nor2_1
X_08693_ _08704_/A _08693_/B VGND VGND VPWR VPWR _08714_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07644_ _07645_/B _07747_/A _07772_/A _07645_/A VGND VGND VPWR VPWR _07646_/A sky130_fd_sc_hd__a22oi_1
XFILLER_54_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07575_ _09215_/A VGND VGND VPWR VPWR _07575_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09314_ _09314_/A VGND VGND VPWR VPWR _12784_/D sky130_fd_sc_hd__clkbuf_1
X_06526_ _06524_/X _06537_/A VGND VGND VPWR VPWR _06529_/A sky130_fd_sc_hd__and2b_1
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09245_ _09195_/A _09242_/X _09244_/Y VGND VGND VPWR VPWR _09256_/A sky130_fd_sc_hd__o21ai_4
X_06457_ _06543_/A _06544_/B _06482_/A VGND VGND VPWR VPWR _06460_/B sky130_fd_sc_hd__a21o_1
X_09176_ _13537_/Q _09183_/B VGND VGND VPWR VPWR _09189_/A sky130_fd_sc_hd__xnor2_1
X_06388_ _12876_/Q VGND VGND VPWR VPWR _10679_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08127_ _14012_/Q _08142_/A VGND VGND VPWR VPWR _08270_/B sky130_fd_sc_hd__and2_1
X_08058_ _12966_/Q _13266_/Q _08062_/S VGND VGND VPWR VPWR _08059_/A sky130_fd_sc_hd__mux2_1
Xoutput36 _13333_/Q VGND VGND VPWR VPWR data_o[15] sky130_fd_sc_hd__buf_2
XFILLER_162_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07009_ hold187/A VGND VGND VPWR VPWR _07063_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput47 _13321_/Q VGND VGND VPWR VPWR data_o[3] sky130_fd_sc_hd__buf_2
XFILLER_103_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10020_ _10020_/A VGND VGND VPWR VPWR _13911_/D sky130_fd_sc_hd__inv_2
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11971_ _11971_/A VGND VGND VPWR VPWR _14300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13710_ _14250_/CLK _13710_/D VGND VGND VPWR VPWR _13710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10922_ _11163_/A VGND VGND VPWR VPWR _10922_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14690_ _14690_/CLK hold442/X VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13641_ _14327_/CLK hold251/X VGND VGND VPWR VPWR _13641_/Q sky130_fd_sc_hd__dfxtp_1
X_10853_ _10853_/A VGND VGND VPWR VPWR _13186_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13572_ _14098_/CLK hold157/X VGND VGND VPWR VPWR _13572_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10784_ _13013_/Q _10790_/B VGND VGND VPWR VPWR _10785_/A sky130_fd_sc_hd__and2_1
XFILLER_9_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12523_ _12545_/A VGND VGND VPWR VPWR _12532_/S sky130_fd_sc_hd__buf_2
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12454_ _12454_/A VGND VGND VPWR VPWR _14658_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11405_ _13726_/Q _11405_/B VGND VGND VPWR VPWR _11406_/A sky130_fd_sc_hd__and2_1
XFILLER_138_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12385_ _12385_/A VGND VGND VPWR VPWR _14614_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14124_ _14716_/CLK hold241/X VGND VGND VPWR VPWR _14124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11336_ _13888_/Q _13885_/Q _11335_/Y VGND VGND VPWR VPWR _12004_/A sky130_fd_sc_hd__a21oi_4
XFILLER_114_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14055_ _14705_/CLK _14055_/D VGND VGND VPWR VPWR _14055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11267_ _11267_/A VGND VGND VPWR VPWR _13390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13006_ _13296_/CLK _13006_/D hold1/X VGND VGND VPWR VPWR _13006_/Q sky130_fd_sc_hd__dfrtp_2
X_10218_ _14098_/Q _14082_/Q _14384_/D VGND VGND VPWR VPWR _10219_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11198_ _11198_/A _11155_/X VGND VGND VPWR VPWR _11198_/X sky130_fd_sc_hd__or2b_1
XFILLER_39_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10149_ _14282_/D _10149_/B VGND VGND VPWR VPWR _10150_/B sky130_fd_sc_hd__nor2_1
XFILLER_82_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13908_ _14210_/CLK _13908_/D VGND VGND VPWR VPWR hold254/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13839_ _14724_/CLK _13839_/D VGND VGND VPWR VPWR _13839_/Q sky130_fd_sc_hd__dfxtp_1
X_07360_ _07343_/X _07358_/Y _07359_/X VGND VGND VPWR VPWR _13138_/D sky130_fd_sc_hd__a21o_1
X_06311_ _13876_/Q _13860_/Q _06313_/S VGND VGND VPWR VPWR _06312_/A sky130_fd_sc_hd__mux2_1
X_07291_ _07305_/A _07290_/X VGND VGND VPWR VPWR _07294_/A sky130_fd_sc_hd__or2b_1
XFILLER_148_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09030_ _09030_/A VGND VGND VPWR VPWR _12751_/D sky130_fd_sc_hd__clkbuf_1
X_06242_ _06242_/A VGND VGND VPWR VPWR _14390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06173_ _13860_/Q _06175_/B VGND VGND VPWR VPWR _06174_/A sky130_fd_sc_hd__and2_1
Xhold302 hold302/A VGND VGND VPWR VPWR hold302/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_117_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold313 hold313/A VGND VGND VPWR VPWR hold313/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold324 hold324/A VGND VGND VPWR VPWR hold324/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold335 hold335/A VGND VGND VPWR VPWR hold335/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold346 hold346/A VGND VGND VPWR VPWR hold346/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold357 hold357/A VGND VGND VPWR VPWR hold357/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_117_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold368 hold368/A VGND VGND VPWR VPWR hold368/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09932_ _09932_/A VGND VGND VPWR VPWR _12853_/D sky130_fd_sc_hd__clkbuf_1
Xhold379 hold379/A VGND VGND VPWR VPWR hold379/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_98_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _13687_/Q _09870_/B VGND VGND VPWR VPWR _09865_/A sky130_fd_sc_hd__and2_1
XFILLER_112_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08814_ _08851_/A _08927_/A _08833_/C VGND VGND VPWR VPWR _08816_/A sky130_fd_sc_hd__and3_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _09781_/Y _09773_/B _09780_/A _09770_/A VGND VGND VPWR VPWR _09795_/B sky130_fd_sc_hd__a211o_1
XFILLER_85_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08745_ _08689_/B _08742_/Y _08744_/X VGND VGND VPWR VPWR _08758_/A sky130_fd_sc_hd__a21o_1
XFILLER_100_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05957_ _13631_/Q _13632_/Q _13633_/Q _13634_/Q VGND VGND VPWR VPWR _05957_/X sky130_fd_sc_hd__and4_1
XFILLER_100_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08676_ _09524_/B VGND VGND VPWR VPWR _09525_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _07701_/B _07723_/A _07627_/C VGND VGND VPWR VPWR _07656_/A sky130_fd_sc_hd__and3_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07558_ _07399_/X _07557_/Y _07475_/X VGND VGND VPWR VPWR _13158_/D sky130_fd_sc_hd__a21o_1
XFILLER_42_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06509_ _06505_/B _06508_/X _06530_/S VGND VGND VPWR VPWR _06510_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07489_ _13149_/Q _07513_/B VGND VGND VPWR VPWR _07498_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09228_ _13544_/Q _09228_/B VGND VGND VPWR VPWR _09228_/X sky130_fd_sc_hd__or2_1
XFILLER_6_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09159_ _09159_/A _09159_/B _09159_/C VGND VGND VPWR VPWR _09160_/B sky130_fd_sc_hd__or3_1
XFILLER_107_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12170_ _14497_/Q _11978_/X _12172_/S VGND VGND VPWR VPWR _12171_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11121_ _11177_/A _11121_/B VGND VGND VPWR VPWR _11121_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11052_ _11108_/A _11052_/B VGND VGND VPWR VPWR _11052_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10003_ _10003_/A VGND VGND VPWR VPWR _12668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14742_ _14742_/CLK _14742_/D VGND VGND VPWR VPWR _14742_/Q sky130_fd_sc_hd__dfxtp_1
X_11954_ _14295_/Q _11950_/X _11966_/S VGND VGND VPWR VPWR _11955_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10905_ _12566_/A VGND VGND VPWR VPWR _11185_/A sky130_fd_sc_hd__buf_2
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14673_ _14688_/CLK _14673_/D VGND VGND VPWR VPWR hold278/A sky130_fd_sc_hd__dfxtp_1
X_11885_ _11885_/A VGND VGND VPWR VPWR _14239_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_192_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _14579_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13624_ _13635_/CLK hold100/X VGND VGND VPWR VPWR _13624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10836_ _10836_/A VGND VGND VPWR VPWR _13178_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13555_ _13555_/CLK _13555_/D repeater57/X VGND VGND VPWR VPWR _13555_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10767_ _10767_/A VGND VGND VPWR VPWR _13047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12506_ _14076_/Q VGND VGND VPWR VPWR _12506_/Y sky130_fd_sc_hd__inv_2
X_13486_ _13721_/CLK hold168/X VGND VGND VPWR VPWR _13486_/Q sky130_fd_sc_hd__dfxtp_1
X_10698_ _12885_/Q _10698_/B VGND VGND VPWR VPWR _10699_/A sky130_fd_sc_hd__and2_1
XFILLER_139_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12437_ _14651_/Q _14697_/Q _12439_/S VGND VGND VPWR VPWR _12438_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12368_ _12368_/A VGND VGND VPWR VPWR _14606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14107_ _14108_/CLK _14107_/D VGND VGND VPWR VPWR _14107_/Q sky130_fd_sc_hd__dfxtp_1
X_11319_ _11319_/A VGND VGND VPWR VPWR _13766_/D sky130_fd_sc_hd__clkbuf_1
X_12299_ _12299_/A VGND VGND VPWR VPWR _14565_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14038_ _14050_/CLK _14038_/D VGND VGND VPWR VPWR _14038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06860_ _06665_/X _06856_/Y _06870_/B _06859_/X VGND VGND VPWR VPWR _13012_/D sky130_fd_sc_hd__a31o_1
XFILLER_94_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06791_ _06791_/A _06826_/A VGND VGND VPWR VPWR _06827_/B sky130_fd_sc_hd__or2_1
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08530_ _08530_/A _08530_/B VGND VGND VPWR VPWR _08531_/B sky130_fd_sc_hd__and2_1
XFILLER_36_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08461_ _08454_/X _08459_/X _09502_/A VGND VGND VPWR VPWR _08462_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_183_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _14742_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07412_ _13141_/Q _09151_/B _07414_/B VGND VGND VPWR VPWR _07412_/X sky130_fd_sc_hd__a21o_1
X_08392_ _08392_/A VGND VGND VPWR VPWR _12728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07343_ _08296_/B VGND VGND VPWR VPWR _07343_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07274_ _09093_/B VGND VGND VPWR VPWR _09101_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09013_ _09013_/A VGND VGND VPWR VPWR _12743_/D sky130_fd_sc_hd__clkbuf_1
X_06225_ _14396_/Q _14388_/Q _10197_/A VGND VGND VPWR VPWR _10626_/B sky130_fd_sc_hd__mux2_1
XFILLER_163_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold110 hold110/A VGND VGND VPWR VPWR hold110/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06156_ _14183_/Q _14175_/Q _06289_/S VGND VGND VPWR VPWR _06156_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold121 hold121/A VGND VGND VPWR VPWR hold121/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold132 hold132/A VGND VGND VPWR VPWR hold132/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold143 hold143/A VGND VGND VPWR VPWR hold143/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_105_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold154 hold154/A VGND VGND VPWR VPWR hold154/X sky130_fd_sc_hd__clkbuf_1
XFILLER_144_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold165 hold165/A VGND VGND VPWR VPWR hold165/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_06087_ _10606_/B _06086_/X _10034_/S VGND VGND VPWR VPWR _06088_/A sky130_fd_sc_hd__mux2_1
Xhold176 hold176/A VGND VGND VPWR VPWR hold176/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold187 hold187/A VGND VGND VPWR VPWR hold187/X sky130_fd_sc_hd__clkbuf_2
Xhold198 hold198/A VGND VGND VPWR VPWR hold198/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_99_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09915_ _09974_/S VGND VGND VPWR VPWR _09924_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_58_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09846_ _09840_/Y _09833_/B _09842_/A _09845_/X VGND VGND VPWR VPWR _09858_/C sky130_fd_sc_hd__a31o_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09777_ _13676_/Q _09778_/C _09809_/C VGND VGND VPWR VPWR _09780_/A sky130_fd_sc_hd__and3_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06989_ _06987_/Y _06988_/X _06930_/X VGND VGND VPWR VPWR _13026_/D sky130_fd_sc_hd__o21bai_1
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _08728_/A _08724_/B VGND VGND VPWR VPWR _08728_/X sky130_fd_sc_hd__or2b_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _09471_/B VGND VGND VPWR VPWR _09472_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_174_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _14539_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11670_ _14018_/Q _11465_/X _11678_/S VGND VGND VPWR VPWR _11671_/A sky130_fd_sc_hd__mux2_1
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10621_ _14288_/Q _14287_/Q VGND VGND VPWR VPWR _10621_/X sky130_fd_sc_hd__or2_1
XFILLER_41_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13340_ _14619_/CLK _13340_/D VGND VGND VPWR VPWR _13340_/Q sky130_fd_sc_hd__dfxtp_4
X_10552_ _10553_/A _10553_/B VGND VGND VPWR VPWR _14436_/D sky130_fd_sc_hd__xor2_1
XFILLER_6_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13271_ _13273_/CLK _13271_/D repeater59/X VGND VGND VPWR VPWR _13271_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_10_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10483_ _10495_/A _10483_/B VGND VGND VPWR VPWR _10485_/C sky130_fd_sc_hd__and2_1
X_12222_ _12220_/X _12222_/B _12222_/C VGND VGND VPWR VPWR _12223_/A sky130_fd_sc_hd__and3b_1
XFILLER_163_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12153_ _14489_/Q _11950_/X _12161_/S VGND VGND VPWR VPWR _12154_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11104_ _11104_/A VGND VGND VPWR VPWR _11104_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12084_ _12084_/A VGND VGND VPWR VPWR _14459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11035_ _11035_/A _11035_/B VGND VGND VPWR VPWR _11035_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12986_ _14633_/CLK hold516/X VGND VGND VPWR VPWR _13107_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_33_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14725_ _14725_/CLK _14725_/D VGND VGND VPWR VPWR _14725_/Q sky130_fd_sc_hd__dfxtp_1
X_11937_ _11937_/A VGND VGND VPWR VPWR _14274_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_165_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _14557_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_150_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11868_ _11868_/A VGND VGND VPWR VPWR _14231_/D sky130_fd_sc_hd__clkbuf_1
X_14656_ _14656_/CLK _14656_/D VGND VGND VPWR VPWR _14656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10819_ _10819_/A VGND VGND VPWR VPWR _13071_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_13607_ _13610_/CLK _13607_/D repeater57/X VGND VGND VPWR VPWR _13607_/Q sky130_fd_sc_hd__dfrtp_2
X_14587_ _14688_/CLK _14587_/D VGND VGND VPWR VPWR hold288/A sky130_fd_sc_hd__dfxtp_1
X_11799_ _11799_/A VGND VGND VPWR VPWR _14092_/D sky130_fd_sc_hd__clkbuf_1
X_13538_ _13558_/CLK _13538_/D _12609_/A VGND VGND VPWR VPWR _13538_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_119_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13469_ _13621_/CLK _13469_/D VGND VGND VPWR VPWR _13469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06010_ _13575_/Q _13580_/Q _13581_/Q _13582_/Q VGND VGND VPWR VPWR _06012_/B sky130_fd_sc_hd__and4_1
XFILLER_127_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07961_ _07948_/A _07952_/X _07957_/B VGND VGND VPWR VPWR _07961_/X sky130_fd_sc_hd__a21bo_1
XFILLER_87_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09700_ _14219_/Q _14217_/Q _09715_/S VGND VGND VPWR VPWR _09700_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06912_ _06919_/A _06912_/B VGND VGND VPWR VPWR _06924_/C sky130_fd_sc_hd__nand2_1
XFILLER_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07892_ _07892_/A _07892_/B _07892_/C _07892_/D VGND VGND VPWR VPWR _07893_/C sky130_fd_sc_hd__or4_1
XFILLER_68_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09631_ _13412_/Q _13610_/Q _09631_/S VGND VGND VPWR VPWR _09632_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06843_ _06843_/A VGND VGND VPWR VPWR _07895_/C sky130_fd_sc_hd__clkbuf_1
X_09562_ _13617_/Q _09562_/B VGND VGND VPWR VPWR _09564_/A sky130_fd_sc_hd__and2_1
XFILLER_83_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06774_ _13006_/Q _06781_/B VGND VGND VPWR VPWR _06827_/A sky130_fd_sc_hd__xnor2_1
X_08513_ _08512_/A _08512_/C _08512_/B VGND VGND VPWR VPWR _08513_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_24_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09493_ _09493_/A VGND VGND VPWR VPWR _09493_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_156_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _14657_/CLK sky130_fd_sc_hd__clkbuf_16
X_08444_ _14252_/Q _14250_/Q _13474_/Q VGND VGND VPWR VPWR _08444_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08375_ _08397_/A VGND VGND VPWR VPWR _08384_/S sky130_fd_sc_hd__buf_2
X_07326_ _07396_/A VGND VGND VPWR VPWR _07326_/X sky130_fd_sc_hd__buf_2
XFILLER_164_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07257_ _07258_/A _07258_/B VGND VGND VPWR VPWR _07257_/X sky130_fd_sc_hd__or2_1
X_06208_ _06208_/A VGND VGND VPWR VPWR _14370_/D sky130_fd_sc_hd__clkbuf_1
X_07188_ _07165_/A _07203_/B _07166_/A _07164_/B VGND VGND VPWR VPWR _07204_/A sky130_fd_sc_hd__a31o_1
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06139_ _14191_/Q _14183_/Q _14194_/D VGND VGND VPWR VPWR _06292_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09829_ _13681_/Q _09829_/B VGND VGND VPWR VPWR _09830_/B sky130_fd_sc_hd__nor2_1
XFILLER_46_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12840_ _14657_/CLK _12840_/D VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__dfxtp_1
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _13698_/CLK _12771_/D VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__dfxtp_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_147_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _14716_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ _14510_/CLK _14510_/D VGND VGND VPWR VPWR _14510_/Q sky130_fd_sc_hd__dfxtp_1
X_11722_ _11722_/A VGND VGND VPWR VPWR _14053_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14441_ _14742_/CLK _14441_/D VGND VGND VPWR VPWR _14441_/Q sky130_fd_sc_hd__dfxtp_1
X_11653_ _14002_/Q _11522_/X _11653_/S VGND VGND VPWR VPWR _11654_/A sky130_fd_sc_hd__mux2_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10604_ _14045_/Q _13914_/Q _13922_/Q _13895_/Q VGND VGND VPWR VPWR _10604_/X sky130_fd_sc_hd__or4_1
X_14372_ _14536_/CLK hold366/X VGND VGND VPWR VPWR hold356/A sky130_fd_sc_hd__dfxtp_1
X_11584_ _11584_/A VGND VGND VPWR VPWR _13873_/D sky130_fd_sc_hd__clkbuf_1
X_13323_ _14712_/CLK _13323_/D VGND VGND VPWR VPWR _13323_/Q sky130_fd_sc_hd__dfxtp_4
X_10535_ _10547_/A _10534_/B _10533_/X VGND VGND VPWR VPWR _10536_/B sky130_fd_sc_hd__o21bai_1
XFILLER_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13254_ _13258_/CLK _13254_/D hold1/X VGND VGND VPWR VPWR _13254_/Q sky130_fd_sc_hd__dfrtp_1
X_10466_ _10466_/A _10466_/B VGND VGND VPWR VPWR _10468_/B sky130_fd_sc_hd__nor2_1
XFILLER_124_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12205_ _12222_/B VGND VGND VPWR VPWR _12205_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13185_ _13423_/CLK _13185_/D VGND VGND VPWR VPWR hold376/A sky130_fd_sc_hd__dfxtp_1
X_10397_ _10397_/A _10396_/X VGND VGND VPWR VPWR _10400_/A sky130_fd_sc_hd__or2b_1
X_12136_ _12136_/A VGND VGND VPWR VPWR _14482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12067_ _12067_/A VGND VGND VPWR VPWR _14451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11018_ _14601_/Q _14563_/Q _14494_/Q _14446_/Q _10969_/X _10970_/X VGND VGND VPWR
+ VPWR _11019_/A sky130_fd_sc_hd__mux4_1
XFILLER_49_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_138_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _14292_/CLK sky130_fd_sc_hd__clkbuf_16
X_12969_ _13273_/CLK hold133/X VGND VGND VPWR VPWR _12969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14708_ _14710_/CLK _14708_/D VGND VGND VPWR VPWR _14708_/Q sky130_fd_sc_hd__dfxtp_1
X_06490_ _06490_/A _06490_/B VGND VGND VPWR VPWR _06490_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14639_ _14643_/CLK _14639_/D VGND VGND VPWR VPWR _14639_/Q sky130_fd_sc_hd__dfxtp_1
X_08160_ _08176_/A _08250_/B _08177_/A VGND VGND VPWR VPWR _08164_/B sky130_fd_sc_hd__a21o_1
X_07111_ _07111_/A _07111_/B VGND VGND VPWR VPWR _07113_/A sky130_fd_sc_hd__nor2_1
X_08091_ _12981_/Q _13281_/Q _08095_/S VGND VGND VPWR VPWR _08092_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07042_ _07141_/B VGND VGND VPWR VPWR _07163_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08993_ _08993_/A _08993_/B _08993_/C VGND VGND VPWR VPWR _08994_/B sky130_fd_sc_hd__and3_1
XFILLER_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07944_ _07944_/A _07944_/B _07949_/D VGND VGND VPWR VPWR _07944_/Y sky130_fd_sc_hd__nand3_1
XFILLER_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07875_ _07811_/X _07881_/B _07874_/Y _06808_/X VGND VGND VPWR VPWR _13262_/D sky130_fd_sc_hd__a31o_1
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09614_ _13404_/Q _13602_/Q _09620_/S VGND VGND VPWR VPWR _09615_/A sky130_fd_sc_hd__mux2_1
X_06826_ _06826_/A _06826_/B _06826_/C VGND VGND VPWR VPWR _06826_/X sky130_fd_sc_hd__or3_1
XFILLER_44_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09545_ _08504_/X _09544_/X _09493_/X VGND VGND VPWR VPWR _13614_/D sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_129_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _13978_/CLK sky130_fd_sc_hd__clkbuf_16
X_06757_ _13005_/Q _06757_/B VGND VGND VPWR VPWR _06759_/A sky130_fd_sc_hd__nor2_1
XFILLER_55_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09476_ _09437_/X _09474_/X _09475_/Y _08665_/X VGND VGND VPWR VPWR _13604_/D sky130_fd_sc_hd__a31o_1
X_06688_ _13347_/Q _13343_/Q _13345_/Q _12672_/Q _06674_/C _06746_/S VGND VGND VPWR
+ VPWR _06688_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08427_ _08427_/A VGND VGND VPWR VPWR _08671_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_8_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08358_ _13077_/Q _13358_/Q _08362_/S VGND VGND VPWR VPWR _08359_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07309_ _07224_/A _07428_/B _07243_/X _07244_/X _07372_/S _07327_/A VGND VGND VPWR
+ VPWR _07311_/C sky130_fd_sc_hd__mux4_1
XFILLER_109_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08289_ _08283_/Y _08276_/B _08285_/A _08288_/X VGND VGND VPWR VPWR _08301_/C sky130_fd_sc_hd__a31o_1
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10320_ _13746_/Q _13106_/Q _10321_/C VGND VGND VPWR VPWR _10322_/A sky130_fd_sc_hd__o21a_1
XFILLER_4_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10251_ _10190_/A _10231_/X _10246_/X VGND VGND VPWR VPWR _10251_/X sky130_fd_sc_hd__a21o_1
XFILLER_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10182_ _10179_/X _14140_/D _10182_/S VGND VGND VPWR VPWR _10183_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13941_ _13964_/CLK _13941_/D VGND VGND VPWR VPWR _13941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13872_ _14656_/CLK _13872_/D VGND VGND VPWR VPWR _13872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12823_ _13653_/CLK _12823_/D VGND VGND VPWR VPWR hold489/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _13704_/CLK _12754_/D VGND VGND VPWR VPWR hold129/A sky130_fd_sc_hd__dfxtp_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _11705_/A VGND VGND VPWR VPWR _14034_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12685_ _13296_/CLK _12685_/D VGND VGND VPWR VPWR hold134/A sky130_fd_sc_hd__dfxtp_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14424_ _14424_/CLK _14424_/D VGND VGND VPWR VPWR _14424_/Q sky130_fd_sc_hd__dfxtp_1
X_11636_ _11636_/A VGND VGND VPWR VPWR _11645_/S sky130_fd_sc_hd__buf_2
XFILLER_30_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11567_ _11567_/A VGND VGND VPWR VPWR _13865_/D sky130_fd_sc_hd__clkbuf_1
X_14355_ _14357_/CLK _14355_/D VGND VGND VPWR VPWR hold439/A sky130_fd_sc_hd__dfxtp_1
XFILLER_156_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10518_ _12992_/D _12989_/D VGND VGND VPWR VPWR _10526_/C sky130_fd_sc_hd__and2_1
X_13306_ _13570_/CLK hold422/X VGND VGND VPWR VPWR _13306_/Q sky130_fd_sc_hd__dfxtp_1
X_14286_ _14294_/CLK _14286_/D VGND VGND VPWR VPWR _14286_/Q sky130_fd_sc_hd__dfxtp_1
X_11498_ _11498_/A VGND VGND VPWR VPWR _11511_/S sky130_fd_sc_hd__buf_2
XFILLER_6_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13237_ _13605_/CLK hold517/X VGND VGND VPWR VPWR _13237_/Q sky130_fd_sc_hd__dfxtp_1
X_10449_ _10449_/A _10456_/C VGND VGND VPWR VPWR _10468_/A sky130_fd_sc_hd__and2_1
X_13168_ _13423_/CLK _13168_/D VGND VGND VPWR VPWR _13168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12119_ _12130_/A VGND VGND VPWR VPWR _12128_/S sky130_fd_sc_hd__buf_2
XFILLER_2_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05990_ _14103_/Q _14104_/Q _14105_/Q _14106_/Q VGND VGND VPWR VPWR _05992_/B sky130_fd_sc_hd__and4_1
X_13099_ _14082_/CLK hold451/X VGND VGND VPWR VPWR _13099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07660_ _07683_/A _07660_/B VGND VGND VPWR VPWR _07661_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06611_ _12903_/Q _06620_/B VGND VGND VPWR VPWR _06613_/A sky130_fd_sc_hd__and2_1
XFILLER_81_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07591_ _14702_/Q VGND VGND VPWR VPWR _07613_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09330_ _13302_/Q _13540_/Q _09332_/S VGND VGND VPWR VPWR _09331_/A sky130_fd_sc_hd__mux2_1
X_06542_ _06599_/A VGND VGND VPWR VPWR _06542_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09261_ _09267_/A _09261_/B _09261_/C VGND VGND VPWR VPWR _09261_/Y sky130_fd_sc_hd__nand3_1
X_06473_ _12882_/Q _06473_/B VGND VGND VPWR VPWR _06474_/B sky130_fd_sc_hd__nor2_1
XFILLER_60_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08212_ _08189_/A _08202_/A _08202_/B VGND VGND VPWR VPWR _08212_/Y sky130_fd_sc_hd__o21bai_1
X_09192_ _13538_/Q _09188_/B _09190_/B _09191_/Y VGND VGND VPWR VPWR _09192_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_119_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08143_ _08143_/A VGND VGND VPWR VPWR _08176_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08074_ _08074_/A VGND VGND VPWR VPWR _12697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07025_ _13706_/Q VGND VGND VPWR VPWR _07139_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_76_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08976_ _08953_/A _08991_/B _08954_/A _08952_/B VGND VGND VPWR VPWR _08992_/A sky130_fd_sc_hd__a31o_1
XFILLER_152_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_07927_ _07925_/A _07949_/A _07923_/A VGND VGND VPWR VPWR _07934_/A sky130_fd_sc_hd__o21a_1
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold69 hold69/A VGND VGND VPWR VPWR hold69/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07858_ _07858_/A _07858_/B _07858_/C _07858_/D VGND VGND VPWR VPWR _07859_/D sky130_fd_sc_hd__nor4_2
XFILLER_44_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06809_ _06665_/X _06820_/B _06806_/Y _06808_/X VGND VGND VPWR VPWR _13008_/D sky130_fd_sc_hd__a31o_1
X_07789_ _07789_/A _07789_/B VGND VGND VPWR VPWR _07790_/B sky130_fd_sc_hd__xnor2_1
XFILLER_25_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09528_ _09519_/A _09523_/X _09534_/C _08733_/X VGND VGND VPWR VPWR _09528_/X sky130_fd_sc_hd__a31o_1
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09459_ _09467_/A _09466_/A VGND VGND VPWR VPWR _09478_/A sky130_fd_sc_hd__nor2_1
X_12470_ _14666_/Q _12010_/A _12472_/S VGND VGND VPWR VPWR _12471_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11421_ _13733_/Q _11427_/B VGND VGND VPWR VPWR _11422_/A sky130_fd_sc_hd__and2_1
XFILLER_137_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14140_ _14292_/CLK _14140_/D VGND VGND VPWR VPWR hold393/A sky130_fd_sc_hd__dfxtp_1
X_11352_ _13890_/Q _11351_/C _13891_/Q VGND VGND VPWR VPWR _11353_/C sky130_fd_sc_hd__a21o_1
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10303_ _14645_/Q _14646_/Q VGND VGND VPWR VPWR hold486/A sky130_fd_sc_hd__xnor2_1
X_14071_ _14617_/CLK _14071_/D VGND VGND VPWR VPWR _14071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11283_ _13755_/Q _11272_/X _11295_/S VGND VGND VPWR VPWR _11284_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13022_ _13570_/CLK _13022_/D repeater59/X VGND VGND VPWR VPWR _13022_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_152_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10234_ _10234_/A VGND VGND VPWR VPWR _10237_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10165_ _10151_/X _10164_/X _14293_/D VGND VGND VPWR VPWR _10165_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10096_ _10096_/A VGND VGND VPWR VPWR _13907_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13924_ _14047_/CLK _13924_/D VGND VGND VPWR VPWR hold69/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13855_ _13855_/CLK _13855_/D VGND VGND VPWR VPWR _13855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12806_ _13587_/CLK _12806_/D VGND VGND VPWR VPWR hold222/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10998_ _10998_/A _10925_/X VGND VGND VPWR VPWR _10998_/X sky130_fd_sc_hd__or2b_1
X_13786_ _13799_/CLK _13786_/D VGND VGND VPWR VPWR _13786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _14333_/CLK _12737_/D VGND VGND VPWR VPWR hold85/A sky130_fd_sc_hd__dfxtp_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12668_ _14633_/CLK _12668_/D VGND VGND VPWR VPWR _12990_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14407_ _14410_/CLK _14407_/D VGND VGND VPWR VPWR _14407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11619_ _13986_/Q _11472_/X _11623_/S VGND VGND VPWR VPWR _11620_/A sky130_fd_sc_hd__mux2_1
X_12599_ _14730_/Q _12619_/B VGND VGND VPWR VPWR _12599_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14338_ _14696_/CLK hold113/X VGND VGND VPWR VPWR _14338_/Q sky130_fd_sc_hd__dfxtp_1
Xhold506 hold506/A VGND VGND VPWR VPWR hold506/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold517 hold517/A VGND VGND VPWR VPWR hold517/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14269_ _14716_/CLK _14269_/D VGND VGND VPWR VPWR _14269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08830_ _08929_/B VGND VGND VPWR VPWR _08951_/A sky130_fd_sc_hd__clkbuf_2
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _08767_/A _08761_/B VGND VGND VPWR VPWR _08770_/A sky130_fd_sc_hd__nand2_1
XFILLER_111_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05973_ _13649_/Q _13650_/Q _13651_/Q _13652_/Q VGND VGND VPWR VPWR _05976_/A sky130_fd_sc_hd__or4_1
XFILLER_85_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07712_ _07735_/A _07712_/B VGND VGND VPWR VPWR _07716_/B sky130_fd_sc_hd__or2_1
XFILLER_66_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08692_ _13452_/Q _09525_/B VGND VGND VPWR VPWR _08693_/B sky130_fd_sc_hd__or2_1
XFILLER_54_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07643_ _07723_/C VGND VGND VPWR VPWR _07772_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07574_ _07571_/Y _07572_/X _07566_/A _07567_/Y VGND VGND VPWR VPWR _07574_/X sky130_fd_sc_hd__a211o_1
XFILLER_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09313_ _13294_/Q _13532_/Q _09321_/S VGND VGND VPWR VPWR _09314_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06525_ _12887_/Q _06525_/B VGND VGND VPWR VPWR _06537_/A sky130_fd_sc_hd__or2_1
XFILLER_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_60_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _13524_/CLK sky130_fd_sc_hd__clkbuf_16
X_09244_ _09244_/A _09244_/B VGND VGND VPWR VPWR _09244_/Y sky130_fd_sc_hd__nor2_1
X_06456_ _12671_/Q _14438_/Q _06469_/A VGND VGND VPWR VPWR _06544_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09175_ _09125_/X _09174_/X _07436_/Y VGND VGND VPWR VPWR _13536_/D sky130_fd_sc_hd__a21o_1
XFILLER_119_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06387_ _06446_/A _06387_/B VGND VGND VPWR VPWR _06391_/A sky130_fd_sc_hd__and2_2
XFILLER_147_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08126_ _14010_/Q _14008_/Q _13424_/Q VGND VGND VPWR VPWR _08126_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08057_ _08057_/A VGND VGND VPWR VPWR _12689_/D sky130_fd_sc_hd__clkbuf_1
Xoutput37 _13334_/Q VGND VGND VPWR VPWR data_o[16] sky130_fd_sc_hd__buf_2
X_07008_ _06945_/X _07006_/X _07007_/Y _06974_/X VGND VGND VPWR VPWR _13029_/D sky130_fd_sc_hd__a31o_1
Xoutput48 _13322_/Q VGND VGND VPWR VPWR data_o[4] sky130_fd_sc_hd__buf_2
XFILLER_131_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08959_ _08934_/B _08959_/B VGND VGND VPWR VPWR _08959_/X sky130_fd_sc_hd__and2b_1
XFILLER_76_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11970_ _14300_/Q _11968_/X _11982_/S VGND VGND VPWR VPWR _11971_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10921_ _11162_/A VGND VGND VPWR VPWR _10921_/X sky130_fd_sc_hd__buf_2
XFILLER_84_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13640_ _13653_/CLK hold149/X VGND VGND VPWR VPWR _13640_/Q sky130_fd_sc_hd__dfxtp_1
X_10852_ _13144_/Q _10852_/B VGND VGND VPWR VPWR _10853_/A sky130_fd_sc_hd__and2_1
XFILLER_32_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ _14319_/CLK hold51/X VGND VGND VPWR VPWR _13571_/Q sky130_fd_sc_hd__dfxtp_1
X_10783_ _10783_/A VGND VGND VPWR VPWR _13054_/D sky130_fd_sc_hd__clkbuf_1
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_51_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _14690_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_157_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12522_ _12522_/A VGND VGND VPWR VPWR _14707_/D sky130_fd_sc_hd__clkbuf_1
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12453_ _14658_/Q _14515_/Q _12461_/S VGND VGND VPWR VPWR _12454_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11404_ _11404_/A VGND VGND VPWR VPWR _13794_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12384_ _14614_/Q _12010_/X _12386_/S VGND VGND VPWR VPWR _12385_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11335_ _13888_/Q _13885_/Q _11353_/B VGND VGND VPWR VPWR _11335_/Y sky130_fd_sc_hd__o21ai_1
X_14123_ _14159_/CLK hold237/X VGND VGND VPWR VPWR _14123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14054_ _14705_/CLK _14054_/D VGND VGND VPWR VPWR _14054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11266_ _11266_/A _11266_/B VGND VGND VPWR VPWR _11267_/A sky130_fd_sc_hd__and2_1
XFILLER_79_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10217_ _10217_/A VGND VGND VPWR VPWR _14396_/D sky130_fd_sc_hd__clkbuf_1
X_13005_ _13296_/CLK _13005_/D hold1/X VGND VGND VPWR VPWR _13005_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11197_ _14031_/Q _13997_/Q _13837_/Q _14549_/Q _11152_/X _11153_/X VGND VGND VPWR
+ VPWR _11198_/A sky130_fd_sc_hd__mux4_1
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10148_ _14150_/Q _10143_/X _10150_/A VGND VGND VPWR VPWR _14285_/D sky130_fd_sc_hd__a21o_1
XFILLER_79_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10079_ _10074_/X _10078_/X _14048_/D VGND VGND VPWR VPWR _10080_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13907_ _14209_/CLK _13907_/D VGND VGND VPWR VPWR hold441/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13838_ _14722_/CLK _13838_/D VGND VGND VPWR VPWR _13838_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13769_ _14717_/CLK _13769_/D VGND VGND VPWR VPWR _13769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_42_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _12885_/CLK sky130_fd_sc_hd__clkbuf_16
X_06310_ _06310_/A VGND VGND VPWR VPWR _14189_/D sky130_fd_sc_hd__clkbuf_1
X_07290_ _09099_/A _09099_/B _13134_/Q VGND VGND VPWR VPWR _07290_/X sky130_fd_sc_hd__or3b_1
XFILLER_148_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06241_ _14091_/Q _06245_/B VGND VGND VPWR VPWR _06242_/A sky130_fd_sc_hd__and2_1
XFILLER_164_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06172_ _06172_/A VGND VGND VPWR VPWR _14173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold303 hold303/A VGND VGND VPWR VPWR hold303/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold314 hold314/A VGND VGND VPWR VPWR hold314/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold325 hold325/A VGND VGND VPWR VPWR hold325/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold336 hold336/A VGND VGND VPWR VPWR hold336/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold347 hold347/A VGND VGND VPWR VPWR hold347/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold358 hold358/A VGND VGND VPWR VPWR hold358/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold369 hold369/A VGND VGND VPWR VPWR hold369/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09931_ _13490_/Q _13679_/Q _09935_/S VGND VGND VPWR VPWR _09932_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _09862_/A VGND VGND VPWR VPWR _13686_/D sky130_fd_sc_hd__clkbuf_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08813_ _13517_/D VGND VGND VPWR VPWR _08927_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09793_ _09793_/A VGND VGND VPWR VPWR _09795_/A sky130_fd_sc_hd__inv_2
XFILLER_133_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05956_ _10137_/S VGND VGND VPWR VPWR _14167_/D sky130_fd_sc_hd__buf_2
XFILLER_73_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08744_ _08744_/A _08744_/B VGND VGND VPWR VPWR _08744_/X sky130_fd_sc_hd__or2_1
XFILLER_26_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _08689_/B _08714_/A VGND VGND VPWR VPWR _08675_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07626_ _07645_/B _07701_/B _07723_/A _07701_/A VGND VGND VPWR VPWR _07626_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_26_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07557_ _07559_/B _07557_/B VGND VGND VPWR VPWR _07557_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_33_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _13273_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06508_ _06508_/A _06508_/B VGND VGND VPWR VPWR _06508_/X sky130_fd_sc_hd__xor2_1
XFILLER_10_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07488_ _07488_/A _07483_/B VGND VGND VPWR VPWR _07493_/B sky130_fd_sc_hd__or2b_1
XFILLER_10_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09227_ _13544_/Q _09228_/B VGND VGND VPWR VPWR _09229_/A sky130_fd_sc_hd__and2_1
X_06439_ _06439_/A VGND VGND VPWR VPWR _12879_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09158_ _09156_/A _09159_/B _09159_/C VGND VGND VPWR VPWR _09158_/X sky130_fd_sc_hd__o21ba_1
XFILLER_107_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08109_ _08143_/A _08162_/B VGND VGND VPWR VPWR _08147_/A sky130_fd_sc_hd__and2b_1
X_09089_ _09089_/A _09089_/B _09089_/C VGND VGND VPWR VPWR _09089_/X sky130_fd_sc_hd__or3_1
XFILLER_107_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11120_ _14269_/Q _14660_/Q _13767_/Q _14715_/Q _11091_/X _11092_/X VGND VGND VPWR
+ VPWR _11121_/B sky130_fd_sc_hd__mux4_1
XFILLER_116_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11051_ _11017_/X _11047_/Y _11050_/Y _11024_/X VGND VGND VPWR VPWR _11052_/B sky130_fd_sc_hd__a211o_1
XFILLER_1_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10002_ _10001_/X _09994_/X _10635_/B VGND VGND VPWR VPWR _10003_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14741_ _14742_/CLK _14741_/D VGND VGND VPWR VPWR _14741_/Q sky130_fd_sc_hd__dfxtp_1
X_11953_ _12026_/S VGND VGND VPWR VPWR _11966_/S sky130_fd_sc_hd__buf_2
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10904_ _14729_/Q _10901_/X _10903_/Y VGND VGND VPWR VPWR _12566_/A sky130_fd_sc_hd__o21a_1
X_14672_ _14688_/CLK _14672_/D VGND VGND VPWR VPWR hold270/A sky130_fd_sc_hd__dfxtp_1
X_11884_ _14239_/Q _11507_/X _11886_/S VGND VGND VPWR VPWR _11885_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13623_ _13635_/CLK hold387/X VGND VGND VPWR VPWR _13623_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_3_0_clk clkbuf_2_3_0_clk/A VGND VGND VPWR VPWR clkbuf_3_7_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_10835_ _13136_/Q _10841_/B VGND VGND VPWR VPWR _10836_/A sky130_fd_sc_hd__and2_1
XFILLER_41_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _13562_/CLK sky130_fd_sc_hd__clkbuf_16
X_13554_ _13554_/CLK _13554_/D _12609_/A VGND VGND VPWR VPWR _13554_/Q sky130_fd_sc_hd__dfrtp_2
Xrepeater56 hold1/A VGND VGND VPWR VPWR repeater56/X sky130_fd_sc_hd__buf_12
X_10766_ _13005_/Q _10768_/B VGND VGND VPWR VPWR _10767_/A sky130_fd_sc_hd__and2_1
XFILLER_146_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12505_ _12504_/Y _14374_/Q _14327_/Q VGND VGND VPWR VPWR hold82/A sky130_fd_sc_hd__a21o_1
XFILLER_40_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10697_ _10697_/A VGND VGND VPWR VPWR _12927_/D sky130_fd_sc_hd__clkbuf_1
X_13485_ _13721_/CLK hold190/X VGND VGND VPWR VPWR _13485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12436_ _12436_/A VGND VGND VPWR VPWR _14650_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12367_ _14606_/Q _11984_/X _12375_/S VGND VGND VPWR VPWR _12368_/A sky130_fd_sc_hd__mux2_1
X_14106_ _14108_/CLK _14106_/D VGND VGND VPWR VPWR _14106_/Q sky130_fd_sc_hd__dfxtp_1
X_11318_ _13766_/Q _11317_/X _11327_/S VGND VGND VPWR VPWR _11319_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12298_ _14565_/Q _11975_/X _12302_/S VGND VGND VPWR VPWR _12299_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14037_ _14050_/CLK hold152/X VGND VGND VPWR VPWR _14037_/Q sky130_fd_sc_hd__dfxtp_1
X_11249_ _11249_/A VGND VGND VPWR VPWR _11249_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06790_ _07863_/B _07863_/C _13007_/Q VGND VGND VPWR VPWR _06826_/A sky130_fd_sc_hd__a21oi_1
XFILLER_67_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08460_ _13469_/Q VGND VGND VPWR VPWR _09502_/A sky130_fd_sc_hd__buf_2
XFILLER_36_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07411_ _08124_/A VGND VGND VPWR VPWR _07411_/X sky130_fd_sc_hd__clkbuf_2
X_08391_ _13092_/Q _13373_/Q _08395_/S VGND VGND VPWR VPWR _08392_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _14410_/CLK sky130_fd_sc_hd__clkbuf_16
X_07342_ _07326_/X _07356_/B _07338_/X _07341_/Y VGND VGND VPWR VPWR _13137_/D sky130_fd_sc_hd__a22o_1
XFILLER_149_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07273_ _13133_/Q _09093_/B VGND VGND VPWR VPWR _07276_/B sky130_fd_sc_hd__nor2_1
X_09012_ _13207_/Q _13436_/Q _09018_/S VGND VGND VPWR VPWR _09013_/A sky130_fd_sc_hd__mux2_1
X_06224_ _06224_/A VGND VGND VPWR VPWR _14415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold100 hold100/A VGND VGND VPWR VPWR hold100/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_163_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06155_ _14179_/Q _14171_/Q _10110_/A VGND VGND VPWR VPWR _10616_/B sky130_fd_sc_hd__mux2_1
Xhold111 hold111/A VGND VGND VPWR VPWR hold111/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold122 hold122/A VGND VGND VPWR VPWR hold122/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold133 hold133/A VGND VGND VPWR VPWR hold133/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold144 hold144/A VGND VGND VPWR VPWR hold144/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_06086_ _13951_/Q _13943_/Q _06256_/S VGND VGND VPWR VPWR _06086_/X sky130_fd_sc_hd__mux2_1
Xhold155 hold155/A VGND VGND VPWR VPWR hold155/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold166 hold166/A VGND VGND VPWR VPWR hold166/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold177 hold177/A VGND VGND VPWR VPWR hold177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 hold188/A VGND VGND VPWR VPWR hold188/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold199 hold199/A VGND VGND VPWR VPWR hold199/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_09914_ _09914_/A VGND VGND VPWR VPWR _12845_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09845_ _09830_/A _09839_/A _09839_/B VGND VGND VPWR VPWR _09845_/X sky130_fd_sc_hd__o21ba_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09776_ _09855_/A VGND VGND VPWR VPWR _09776_/X sky130_fd_sc_hd__buf_2
XFILLER_160_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06988_ _06996_/A _06996_/B _06836_/X VGND VGND VPWR VPWR _06988_/X sky130_fd_sc_hd__a21o_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ _08706_/X _08725_/X _08726_/Y _08696_/X VGND VGND VPWR VPWR _13456_/D sky130_fd_sc_hd__a31o_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05939_ _11382_/B VGND VGND VPWR VPWR _13931_/D sky130_fd_sc_hd__inv_2
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _09424_/B _08596_/B _08607_/C _08657_/X _08566_/B VGND VGND VPWR VPWR _09471_/B
+ sky130_fd_sc_hd__o311a_2
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _07622_/A _07721_/A _07627_/C VGND VGND VPWR VPWR _07610_/B sky130_fd_sc_hd__a21oi_1
XFILLER_14_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08589_ _08633_/A _08589_/B VGND VGND VPWR VPWR _08589_/Y sky130_fd_sc_hd__nand2_1
X_10620_ _14284_/Q _14283_/Q _14286_/Q _14285_/Q VGND VGND VPWR VPWR _10620_/X sky130_fd_sc_hd__or4_1
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10551_ _10539_/X _10542_/B _10540_/A VGND VGND VPWR VPWR _10553_/B sky130_fd_sc_hd__a21oi_1
XFILLER_50_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10482_ _10485_/B VGND VGND VPWR VPWR _10501_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13270_ _13273_/CLK _13270_/D repeater59/X VGND VGND VPWR VPWR _13270_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12221_ _14124_/Q _12220_/C _14125_/Q VGND VGND VPWR VPWR _12222_/C sky130_fd_sc_hd__a21o_1
XFILLER_163_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12152_ _12202_/S VGND VGND VPWR VPWR _12161_/S sky130_fd_sc_hd__buf_2
XFILLER_2_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11103_ _14607_/Q _14569_/Q _14500_/Q _14452_/Q _11044_/X _11045_/X VGND VGND VPWR
+ VPWR _11104_/A sky130_fd_sc_hd__mux4_1
XFILLER_1_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12083_ _11348_/X _14459_/Q _12085_/S VGND VGND VPWR VPWR _12084_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11034_ _14263_/Q _14654_/Q _13761_/Q _14709_/Q _11020_/X _11021_/X VGND VGND VPWR
+ VPWR _11035_/B sky130_fd_sc_hd__mux4_1
XFILLER_49_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12985_ _14633_/CLK hold203/X VGND VGND VPWR VPWR _13106_/D sky130_fd_sc_hd__dfxtp_2
X_14724_ _14724_/CLK _14724_/D VGND VGND VPWR VPWR _14724_/Q sky130_fd_sc_hd__dfxtp_1
X_11936_ _14274_/Q _11504_/X _11940_/S VGND VGND VPWR VPWR _11937_/A sky130_fd_sc_hd__mux2_1
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14655_ _14710_/CLK _14655_/D VGND VGND VPWR VPWR _14655_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11867_ _14231_/Q _11481_/X _11875_/S VGND VGND VPWR VPWR _11868_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13606_ _13606_/CLK _13606_/D repeater57/X VGND VGND VPWR VPWR _13606_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_159_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10818_ _13029_/Q _10818_/B VGND VGND VPWR VPWR _10819_/A sky130_fd_sc_hd__and2_1
X_14586_ _14688_/CLK hold288/X VGND VGND VPWR VPWR hold519/A sky130_fd_sc_hd__dfxtp_2
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11798_ _13570_/Q _11806_/B VGND VGND VPWR VPWR _11799_/A sky130_fd_sc_hd__and2_1
X_13537_ _13554_/CLK _13537_/D _12609_/A VGND VGND VPWR VPWR _13537_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_119_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10749_ _10749_/A VGND VGND VPWR VPWR _12951_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13468_ _13562_/CLK _13468_/D VGND VGND VPWR VPWR _13700_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12419_ _12419_/A VGND VGND VPWR VPWR _14643_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13399_ _13596_/CLK hold455/X VGND VGND VPWR VPWR _13399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07960_ _07958_/X _07959_/Y _07932_/X VGND VGND VPWR VPWR _13273_/D sky130_fd_sc_hd__a21o_1
XFILLER_114_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _14720_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06911_ _13016_/Q _07963_/B VGND VGND VPWR VPWR _06912_/B sky130_fd_sc_hd__or2_1
X_07891_ _07893_/B _07884_/X _07887_/Y _07893_/A VGND VGND VPWR VPWR _07898_/B sky130_fd_sc_hd__a31o_1
XFILLER_110_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09630_ _09630_/A VGND VGND VPWR VPWR _12828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06842_ _06747_/Y _06841_/Y _06745_/X VGND VGND VPWR VPWR _06843_/A sky130_fd_sc_hd__o21ai_2
XFILLER_110_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09561_ _09548_/A _09548_/B _09559_/Y _09560_/X VGND VGND VPWR VPWR _09574_/A sky130_fd_sc_hd__a31oi_2
X_06773_ _06773_/A VGND VGND VPWR VPWR _06781_/B sky130_fd_sc_hd__clkbuf_2
X_08512_ _08512_/A _08512_/B _08512_/C VGND VGND VPWR VPWR _08530_/B sky130_fd_sc_hd__or3_1
XFILLER_51_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09492_ _09495_/A _09509_/B VGND VGND VPWR VPWR _09492_/X sky130_fd_sc_hd__xor2_1
XFILLER_23_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08443_ _14256_/Q _14254_/Q _13474_/Q VGND VGND VPWR VPWR _08635_/B sky130_fd_sc_hd__mux2_1
XFILLER_149_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08374_ _08374_/A VGND VGND VPWR VPWR _12720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07325_ _07473_/A VGND VGND VPWR VPWR _07396_/A sky130_fd_sc_hd__buf_2
XFILLER_109_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07256_ _13131_/Q _09088_/B VGND VGND VPWR VPWR _07258_/B sky130_fd_sc_hd__nand2_1
X_06207_ _06206_/X _06203_/X _10193_/A VGND VGND VPWR VPWR _06208_/A sky130_fd_sc_hd__mux2_1
X_07187_ _07182_/A _07182_/B _07182_/C VGND VGND VPWR VPWR _07196_/B sky130_fd_sc_hd__a21o_1
XFILLER_152_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06138_ _06138_/A VGND VGND VPWR VPWR _14153_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06069_ _13959_/Q _13951_/Q _13962_/D VGND VGND VPWR VPWR _06259_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09828_ _13681_/Q _09829_/B VGND VGND VPWR VPWR _09830_/A sky130_fd_sc_hd__and2_1
XFILLER_100_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09759_ _13674_/Q _09760_/B VGND VGND VPWR VPWR _09761_/A sky130_fd_sc_hd__and2_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _13698_/CLK _12770_/D VGND VGND VPWR VPWR hold397/A sky130_fd_sc_hd__dfxtp_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _11288_/X _14053_/Q _11725_/S VGND VGND VPWR VPWR _11722_/A sky130_fd_sc_hd__mux2_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _14440_/CLK _14440_/D VGND VGND VPWR VPWR _14440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11652_ _11652_/A VGND VGND VPWR VPWR _14001_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10603_ _14037_/Q _14047_/Q VGND VGND VPWR VPWR _10603_/X sky130_fd_sc_hd__and2_1
X_14371_ _14536_/CLK hold356/X VGND VGND VPWR VPWR _14371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11583_ _13649_/Q _11585_/B VGND VGND VPWR VPWR _11584_/A sky130_fd_sc_hd__and2_1
XFILLER_156_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13322_ _14742_/CLK _13322_/D VGND VGND VPWR VPWR _13322_/Q sky130_fd_sc_hd__dfxtp_4
X_10534_ _10547_/A _10534_/B _10533_/X VGND VGND VPWR VPWR _10549_/A sky130_fd_sc_hd__or3b_1
XFILLER_6_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10465_ _10465_/A _10465_/B VGND VGND VPWR VPWR _10466_/B sky130_fd_sc_hd__nor2_1
XFILLER_6_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13253_ _14690_/CLK _13253_/D hold1/X VGND VGND VPWR VPWR _13253_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12204_ _14076_/Q _14110_/Q VGND VGND VPWR VPWR _12222_/B sky130_fd_sc_hd__nor2_1
X_10396_ _10396_/A _10411_/A VGND VGND VPWR VPWR _10396_/X sky130_fd_sc_hd__or2_1
X_13184_ _13423_/CLK _13184_/D VGND VGND VPWR VPWR hold518/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12135_ _14482_/Q _12007_/X _12139_/S VGND VGND VPWR VPWR _12136_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12066_ _11313_/X _14451_/Q _12074_/S VGND VGND VPWR VPWR _12067_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11017_ _11207_/A VGND VGND VPWR VPWR _11017_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12968_ _12970_/CLK hold359/X VGND VGND VPWR VPWR _12968_/Q sky130_fd_sc_hd__dfxtp_1
X_14707_ _14707_/CLK _14707_/D VGND VGND VPWR VPWR _14707_/Q sky130_fd_sc_hd__dfxtp_1
X_11919_ _11919_/A VGND VGND VPWR VPWR _14266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12899_ _12974_/CLK _12899_/D hold1/X VGND VGND VPWR VPWR _12899_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14638_ _14647_/CLK _14638_/D VGND VGND VPWR VPWR _14638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14569_ _14714_/CLK _14569_/D VGND VGND VPWR VPWR _14569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07110_ hold515/A _13112_/D _07141_/C _14630_/Q VGND VGND VPWR VPWR _07111_/B sky130_fd_sc_hd__and4_1
X_08090_ _08090_/A VGND VGND VPWR VPWR _12704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07041_ hold177/A VGND VGND VPWR VPWR _07141_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08992_ _08992_/A _08992_/B VGND VGND VPWR VPWR _08994_/A sky130_fd_sc_hd__and2_1
XFILLER_88_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07943_ _07944_/A _07944_/B _07949_/D VGND VGND VPWR VPWR _07943_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07874_ _07892_/A _07892_/C _07892_/B VGND VGND VPWR VPWR _07874_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09613_ _09613_/A VGND VGND VPWR VPWR _12820_/D sky130_fd_sc_hd__clkbuf_1
X_06825_ _06825_/A _06825_/B _06825_/C VGND VGND VPWR VPWR _06826_/C sky130_fd_sc_hd__or3_1
XFILLER_83_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09544_ _09547_/B _09544_/B VGND VGND VPWR VPWR _09544_/X sky130_fd_sc_hd__xor2_1
XFILLER_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06756_ _07846_/B _07846_/C VGND VGND VPWR VPWR _06757_/B sky130_fd_sc_hd__and2_1
XFILLER_37_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09475_ _09475_/A _09475_/B _09477_/B VGND VGND VPWR VPWR _09475_/Y sky130_fd_sc_hd__nand3_1
X_06687_ _13036_/Q _13351_/Q _13353_/Q _13349_/Q _06674_/C _06746_/S VGND VGND VPWR
+ VPWR _06812_/B sky130_fd_sc_hd__mux4_2
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08426_ _13473_/Q VGND VGND VPWR VPWR _08427_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08357_ _08357_/A VGND VGND VPWR VPWR _12712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07308_ _07239_/X _07321_/B _07306_/Y _07307_/X VGND VGND VPWR VPWR _13135_/D sky130_fd_sc_hd__a31o_1
XFILLER_20_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08288_ _08273_/A _08282_/A _08282_/B VGND VGND VPWR VPWR _08288_/X sky130_fd_sc_hd__o21ba_1
XFILLER_4_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07239_ _08296_/B VGND VGND VPWR VPWR _07239_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10250_ _10250_/A VGND VGND VPWR VPWR _14336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10181_ _10181_/A VGND VGND VPWR VPWR _14138_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13940_ _13963_/CLK _13940_/D VGND VGND VPWR VPWR _13940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13871_ _14656_/CLK _13871_/D VGND VGND VPWR VPWR _13871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12822_ _13653_/CLK _12822_/D VGND VGND VPWR VPWR hold421/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ _13722_/CLK _12753_/D VGND VGND VPWR VPWR hold315/A sky130_fd_sc_hd__dfxtp_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _14034_/Q _11516_/X _11708_/S VGND VGND VPWR VPWR _11705_/A sky130_fd_sc_hd__mux2_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _13294_/CLK _12684_/D VGND VGND VPWR VPWR hold248/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _14732_/CLK _14423_/D VGND VGND VPWR VPWR _14423_/Q sky130_fd_sc_hd__dfxtp_1
X_11635_ _11635_/A VGND VGND VPWR VPWR _13993_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14354_ _14357_/CLK _14354_/D VGND VGND VPWR VPWR hold373/A sky130_fd_sc_hd__dfxtp_1
X_11566_ _13641_/Q _11574_/B VGND VGND VPWR VPWR _11567_/A sky130_fd_sc_hd__and2_1
X_13305_ _13570_/CLK hold73/X VGND VGND VPWR VPWR _13305_/Q sky130_fd_sc_hd__dfxtp_1
X_10517_ _10512_/A _10567_/A _10510_/B _10555_/B VGND VGND VPWR VPWR _10520_/A sky130_fd_sc_hd__o2bb2a_1
X_14285_ _14294_/CLK _14285_/D VGND VGND VPWR VPWR _14285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11497_ _14693_/Q VGND VGND VPWR VPWR _11497_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13236_ _13605_/CLK hold201/X VGND VGND VPWR VPWR _13236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10448_ hold64/A hold186/A VGND VGND VPWR VPWR _10456_/C sky130_fd_sc_hd__and2_1
XFILLER_108_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13167_ _13524_/CLK _13167_/D VGND VGND VPWR VPWR _13167_/Q sky130_fd_sc_hd__dfxtp_1
X_10379_ _10376_/A _10376_/C _10378_/X VGND VGND VPWR VPWR _10380_/B sky130_fd_sc_hd__a21o_1
XFILLER_97_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12118_ _12118_/A VGND VGND VPWR VPWR _14474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13098_ _14082_/CLK hold372/X VGND VGND VPWR VPWR _13098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12049_ _12049_/A VGND VGND VPWR VPWR _14443_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06610_ _06610_/A VGND VGND VPWR VPWR _12902_/D sky130_fd_sc_hd__clkbuf_1
X_07590_ _07570_/X _07588_/X _07589_/Y _07575_/X VGND VGND VPWR VPWR _13162_/D sky130_fd_sc_hd__a31o_1
XFILLER_80_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06541_ _06541_/A VGND VGND VPWR VPWR _12888_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09260_ _09261_/B _09261_/C _09267_/A VGND VGND VPWR VPWR _09264_/B sky130_fd_sc_hd__a21o_1
X_06472_ _12882_/Q _06473_/B VGND VGND VPWR VPWR _06493_/A sky130_fd_sc_hd__and2_1
XFILLER_61_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08211_ _08211_/A _08211_/B VGND VGND VPWR VPWR _08223_/A sky130_fd_sc_hd__or2_1
X_09191_ _09173_/A _09172_/B _09177_/X VGND VGND VPWR VPWR _09191_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_147_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08142_ _08142_/A VGND VGND VPWR VPWR _08197_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08073_ _12973_/Q _13273_/Q _08073_/S VGND VGND VPWR VPWR _08074_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07024_ _07024_/A VGND VGND VPWR VPWR _13342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08975_ _08970_/A _08970_/B _08970_/C VGND VGND VPWR VPWR _08984_/B sky130_fd_sc_hd__a21o_1
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_69_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07926_ _07909_/X _07924_/X _07925_/Y _06974_/X VGND VGND VPWR VPWR _13268_/D sky130_fd_sc_hd__a31o_1
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07857_ _07835_/A _07839_/Y _07840_/Y _07858_/C _07858_/D VGND VGND VPWR VPWR _07859_/C
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06808_ _06871_/A _07876_/B VGND VGND VPWR VPWR _06808_/X sky130_fd_sc_hd__and2_1
X_07788_ _07788_/A _07788_/B VGND VGND VPWR VPWR _07789_/B sky130_fd_sc_hd__nor2_1
XFILLER_72_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09527_ _09519_/A _09523_/X _09534_/C VGND VGND VPWR VPWR _09532_/B sky130_fd_sc_hd__a21oi_1
X_06739_ _13004_/Q _07838_/B VGND VGND VPWR VPWR _06739_/Y sky130_fd_sc_hd__xnor2_1
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09458_ _09457_/B _09457_/C _13602_/Q VGND VGND VPWR VPWR _09466_/A sky130_fd_sc_hd__a21oi_1
XFILLER_157_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08409_ _09323_/A VGND VGND VPWR VPWR _08418_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_8_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09389_ _13593_/Q _09394_/B VGND VGND VPWR VPWR _09391_/B sky130_fd_sc_hd__xnor2_1
X_11420_ _11420_/A VGND VGND VPWR VPWR _13801_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11351_ _13890_/Q _13891_/Q _11351_/C VGND VGND VPWR VPWR _11362_/C sky130_fd_sc_hd__and3_2
XFILLER_153_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10302_ _10302_/A VGND VGND VPWR VPWR _13751_/D sky130_fd_sc_hd__clkbuf_1
X_14070_ _14510_/CLK _14070_/D VGND VGND VPWR VPWR _14070_/Q sky130_fd_sc_hd__dfxtp_1
X_11282_ _11376_/S VGND VGND VPWR VPWR _11295_/S sky130_fd_sc_hd__buf_2
XFILLER_152_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13021_ _13031_/CLK _13021_/D repeater59/X VGND VGND VPWR VPWR _13021_/Q sky130_fd_sc_hd__dfrtp_1
X_10233_ _10233_/A VGND VGND VPWR VPWR _14526_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10164_ _10103_/A _10144_/X _10159_/X VGND VGND VPWR VPWR _10164_/X sky130_fd_sc_hd__a21o_1
XFILLER_120_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10095_ _10092_/X _13908_/D _10095_/S VGND VGND VPWR VPWR _10096_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13923_ _14050_/CLK hold69/X VGND VGND VPWR VPWR hold213/A sky130_fd_sc_hd__dfxtp_1
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13854_ _14180_/CLK _13854_/D VGND VGND VPWR VPWR _13854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12805_ _14108_/CLK _12805_/D VGND VGND VPWR VPWR hold249/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13785_ _13945_/CLK _13785_/D VGND VGND VPWR VPWR _13785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10997_ _14017_/Q _13983_/Q _13823_/Q _14535_/Q _10921_/X _10922_/X VGND VGND VPWR
+ VPWR _10998_/A sky130_fd_sc_hd__mux4_1
XFILLER_90_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _14696_/CLK _12736_/D VGND VGND VPWR VPWR hold104/A sky130_fd_sc_hd__dfxtp_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12667_ _13351_/CLK _12667_/D VGND VGND VPWR VPWR _12989_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14406_ _14410_/CLK _14406_/D VGND VGND VPWR VPWR _14406_/Q sky130_fd_sc_hd__dfxtp_1
X_11618_ _11618_/A VGND VGND VPWR VPWR _13985_/D sky130_fd_sc_hd__clkbuf_1
X_12598_ _14730_/Q _12623_/B VGND VGND VPWR VPWR _12604_/C sky130_fd_sc_hd__and2_1
XFILLER_117_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14337_ _14697_/CLK hold17/X VGND VGND VPWR VPWR _14337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11549_ _11549_/A VGND VGND VPWR VPWR _13857_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold507 hold507/A VGND VGND VPWR VPWR hold507/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_143_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold518 hold518/A VGND VGND VPWR VPWR hold518/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_14268_ _14717_/CLK _14268_/D VGND VGND VPWR VPWR _14268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13219_ _13423_/CLK hold358/X VGND VGND VPWR VPWR _13219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14199_ _14210_/CLK _14199_/D VGND VGND VPWR VPWR _14199_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08760_ _13461_/Q _09542_/B VGND VGND VPWR VPWR _08761_/B sky130_fd_sc_hd__or2_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05972_ _14075_/D _13622_/Q _13623_/Q _13624_/Q VGND VGND VPWR VPWR _05977_/B sky130_fd_sc_hd__or4_1
X_07711_ _07733_/B _07710_/B _07710_/C VGND VGND VPWR VPWR _07712_/B sky130_fd_sc_hd__a21oi_1
X_08691_ _13452_/Q _08730_/B VGND VGND VPWR VPWR _08704_/A sky130_fd_sc_hd__nand2_1
XFILLER_54_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07642_ _13247_/D VGND VGND VPWR VPWR _07723_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07573_ _07566_/A _07567_/Y _07571_/Y _07572_/X VGND VGND VPWR VPWR _07573_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_22_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09312_ _09323_/A VGND VGND VPWR VPWR _09321_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_80_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06524_ _12887_/Q _06563_/B _06524_/C VGND VGND VPWR VPWR _06524_/X sky130_fd_sc_hd__and3_1
XFILLER_21_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09243_ _13543_/Q _13544_/Q _13545_/Q _13546_/Q _09250_/B VGND VGND VPWR VPWR _09244_/B
+ sky130_fd_sc_hd__o41a_1
XFILLER_21_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06455_ _06455_/A VGND VGND VPWR VPWR _06543_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09174_ _09190_/A _09174_/B VGND VGND VPWR VPWR _09174_/X sky130_fd_sc_hd__xor2_1
X_06386_ _06392_/A _06495_/C _06382_/X _06429_/B VGND VGND VPWR VPWR _06387_/B sky130_fd_sc_hd__a22o_1
XFILLER_108_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08125_ _07326_/X _08220_/B _08120_/C _08124_/X VGND VGND VPWR VPWR _13355_/D sky130_fd_sc_hd__a31o_1
XFILLER_147_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08056_ _12965_/Q _13265_/Q _08062_/S VGND VGND VPWR VPWR _08057_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07007_ _06999_/A _07005_/Y _07003_/Y _07004_/X VGND VGND VPWR VPWR _07007_/Y sky130_fd_sc_hd__o211ai_1
Xoutput38 _13335_/Q VGND VGND VPWR VPWR data_o[17] sky130_fd_sc_hd__buf_2
Xoutput49 _13323_/Q VGND VGND VPWR VPWR data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_163_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08958_ _08978_/D VGND VGND VPWR VPWR _08991_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07909_ _07909_/A VGND VGND VPWR VPWR _07909_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08889_ _08889_/A _08889_/B VGND VGND VPWR VPWR _08890_/B sky130_fd_sc_hd__xnor2_1
XFILLER_91_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10920_ _14745_/Q VGND VGND VPWR VPWR _11162_/A sky130_fd_sc_hd__buf_6
XFILLER_56_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10851_ _10851_/A VGND VGND VPWR VPWR _13185_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13570_ _13570_/CLK hold402/X VGND VGND VPWR VPWR _13570_/Q sky130_fd_sc_hd__dfxtp_1
X_10782_ _13012_/Q _10790_/B VGND VGND VPWR VPWR _10783_/A sky130_fd_sc_hd__and2_1
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12521_ _11294_/X _14707_/Q _12521_/S VGND VGND VPWR VPWR _12522_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12452_ _12463_/A VGND VGND VPWR VPWR _12461_/S sky130_fd_sc_hd__buf_2
XFILLER_138_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11403_ _13725_/Q _11405_/B VGND VGND VPWR VPWR _11404_/A sky130_fd_sc_hd__and2_1
XFILLER_153_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12383_ _12383_/A VGND VGND VPWR VPWR _14613_/D sky130_fd_sc_hd__clkbuf_1
X_14122_ _14292_/CLK hold301/X VGND VGND VPWR VPWR _14122_/Q sky130_fd_sc_hd__dfxtp_1
X_11334_ _11364_/B VGND VGND VPWR VPWR _11353_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14053_ _14742_/CLK _14053_/D VGND VGND VPWR VPWR _14053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11265_ _13341_/Q _10962_/A _11258_/X _11264_/Y VGND VGND VPWR VPWR _13341_/D sky130_fd_sc_hd__o22a_1
XFILLER_106_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13004_ _13256_/CLK _13004_/D hold1/X VGND VGND VPWR VPWR _13004_/Q sky130_fd_sc_hd__dfrtp_1
X_10216_ _14097_/Q _14081_/Q _14384_/D VGND VGND VPWR VPWR _10217_/A sky130_fd_sc_hd__mux2_1
X_11196_ _14313_/Q _14483_/Q _14239_/Q _14069_/Q _11137_/X _11138_/X VGND VGND VPWR
+ VPWR _11196_/X sky130_fd_sc_hd__mux4_1
X_10147_ _10147_/A VGND VGND VPWR VPWR _10150_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10078_ _10064_/X _10077_/X _14049_/D VGND VGND VPWR VPWR _10078_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13906_ _14693_/CLK _13906_/D VGND VGND VPWR VPWR hold273/A sky130_fd_sc_hd__dfxtp_1
XFILLER_63_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13837_ _14721_/CLK _13837_/D VGND VGND VPWR VPWR _13837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13768_ _14716_/CLK _13768_/D VGND VGND VPWR VPWR _13768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12719_ _13596_/CLK _12719_/D VGND VGND VPWR VPWR hold460/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13699_ _13722_/CLK _13699_/D repeater56/X VGND VGND VPWR VPWR _13699_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06240_ _06240_/A VGND VGND VPWR VPWR _14389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06171_ _13859_/Q _06175_/B VGND VGND VPWR VPWR _06172_/A sky130_fd_sc_hd__and2_1
XFILLER_156_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold304 hold304/A VGND VGND VPWR VPWR hold304/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold315 hold315/A VGND VGND VPWR VPWR hold315/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold326 hold326/A VGND VGND VPWR VPWR hold326/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_117_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold337 hold337/A VGND VGND VPWR VPWR hold337/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold348 hold348/A VGND VGND VPWR VPWR hold348/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_09930_ _09930_/A VGND VGND VPWR VPWR _12852_/D sky130_fd_sc_hd__clkbuf_1
Xhold359 hold359/A VGND VGND VPWR VPWR hold359/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_125_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _09870_/B _09894_/A _09861_/C VGND VGND VPWR VPWR _09862_/A sky130_fd_sc_hd__and3b_1
XFILLER_113_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08812_ _08812_/A VGND VGND VPWR VPWR _14245_/D sky130_fd_sc_hd__clkbuf_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _09792_/A _09804_/A VGND VGND VPWR VPWR _09796_/A sky130_fd_sc_hd__or2_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _13455_/Q _13456_/Q _13457_/Q _13458_/Q _09550_/B VGND VGND VPWR VPWR _08744_/B
+ sky130_fd_sc_hd__o41a_1
X_05955_ _06313_/S VGND VGND VPWR VPWR _10137_/S sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _13451_/Q _08730_/B VGND VGND VPWR VPWR _08714_/A sky130_fd_sc_hd__xnor2_1
XFILLER_54_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07625_ _13245_/D VGND VGND VPWR VPWR _07701_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07556_ _07556_/A _07556_/B VGND VGND VPWR VPWR _07557_/B sky130_fd_sc_hd__nand2_1
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06507_ _12884_/Q _06500_/B _06499_/Y VGND VGND VPWR VPWR _06508_/B sky130_fd_sc_hd__a21oi_1
XFILLER_139_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07487_ _07411_/X _07484_/X _07485_/Y _07486_/X VGND VGND VPWR VPWR _13148_/D sky130_fd_sc_hd__a31o_1
XFILLER_158_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09226_ _09226_/A _09226_/B VGND VGND VPWR VPWR _09230_/A sky130_fd_sc_hd__or2_1
X_06438_ _06450_/B _06437_/X _06622_/B VGND VGND VPWR VPWR _06439_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09157_ _09106_/X _09155_/X _09156_/Y _07409_/X VGND VGND VPWR VPWR _13534_/D sky130_fd_sc_hd__a31o_1
X_06369_ _06044_/B _06371_/B input21/X VGND VGND VPWR VPWR _06369_/X sky130_fd_sc_hd__and3b_1
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08108_ _14004_/Q _14003_/Q _08142_/A VGND VGND VPWR VPWR _08108_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09088_ _13523_/Q _09088_/B VGND VGND VPWR VPWR _09089_/C sky130_fd_sc_hd__nand2_1
XFILLER_123_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08039_ _08039_/A VGND VGND VPWR VPWR _12681_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11050_ _11106_/A _11050_/B VGND VGND VPWR VPWR _11050_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10001_ _14627_/Q _14625_/Q _10636_/A VGND VGND VPWR VPWR _10001_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14740_ _14742_/CLK _14740_/D VGND VGND VPWR VPWR _14740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11952_ _12001_/A VGND VGND VPWR VPWR _12026_/S sky130_fd_sc_hd__buf_2
XFILLER_85_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10903_ _12596_/B _14727_/Q _14729_/Q VGND VGND VPWR VPWR _10903_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14671_ _14726_/CLK _14671_/D VGND VGND VPWR VPWR _14671_/Q sky130_fd_sc_hd__dfxtp_1
X_11883_ _11883_/A VGND VGND VPWR VPWR _14238_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13622_ _13622_/CLK hold329/X VGND VGND VPWR VPWR _13622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10834_ _10834_/A VGND VGND VPWR VPWR _13177_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13553_ _13554_/CLK _13553_/D _12609_/A VGND VGND VPWR VPWR _13553_/Q sky130_fd_sc_hd__dfrtp_4
X_10765_ _10765_/A VGND VGND VPWR VPWR _13046_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater57 _12609_/A VGND VGND VPWR VPWR repeater57/X sky130_fd_sc_hd__buf_12
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12504_ _14320_/Q VGND VGND VPWR VPWR _12504_/Y sky130_fd_sc_hd__inv_2
X_13484_ _13721_/CLK hold171/X VGND VGND VPWR VPWR _13484_/Q sky130_fd_sc_hd__dfxtp_1
X_10696_ _12884_/Q _10698_/B VGND VGND VPWR VPWR _10697_/A sky130_fd_sc_hd__and2_1
XFILLER_157_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12435_ _14650_/Q _14696_/Q _12439_/S VGND VGND VPWR VPWR _12436_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12366_ _12377_/A VGND VGND VPWR VPWR _12375_/S sky130_fd_sc_hd__buf_2
XFILLER_5_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14105_ _14108_/CLK _14105_/D VGND VGND VPWR VPWR _14105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11317_ _14516_/Q VGND VGND VPWR VPWR _11317_/X sky130_fd_sc_hd__clkbuf_2
X_12297_ _12297_/A VGND VGND VPWR VPWR _14564_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14036_ _14725_/CLK _14036_/D VGND VGND VPWR VPWR _14036_/Q sky130_fd_sc_hd__dfxtp_1
X_11248_ _14618_/Q _14580_/Q _14511_/Q _14463_/Q _12586_/A _11092_/A VGND VGND VPWR
+ VPWR _11249_/A sky130_fd_sc_hd__mux4_1
XFILLER_68_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11179_ _11179_/A _11179_/B VGND VGND VPWR VPWR _11179_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07410_ _07399_/X _07408_/Y _07409_/X VGND VGND VPWR VPWR _13142_/D sky130_fd_sc_hd__a21o_1
X_08390_ _08390_/A VGND VGND VPWR VPWR _12727_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07341_ _07341_/A _07341_/B VGND VGND VPWR VPWR _07341_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07272_ _09086_/B _07284_/B VGND VGND VPWR VPWR _09093_/B sky130_fd_sc_hd__xor2_2
XFILLER_164_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09011_ _09011_/A VGND VGND VPWR VPWR _12742_/D sky130_fd_sc_hd__clkbuf_1
X_06223_ _10626_/A _06222_/X _10208_/S VGND VGND VPWR VPWR _06224_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06154_ _06154_/A VGND VGND VPWR VPWR _14198_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold101 hold101/A VGND VGND VPWR VPWR hold101/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold112 hold112/A VGND VGND VPWR VPWR hold112/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_117_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold123 hold123/A VGND VGND VPWR VPWR hold123/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold134 hold134/A VGND VGND VPWR VPWR hold134/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06085_ _13947_/Q _13939_/Q _10023_/A VGND VGND VPWR VPWR _10606_/B sky130_fd_sc_hd__mux2_1
Xhold145 hold145/A VGND VGND VPWR VPWR hold145/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold156 hold156/A VGND VGND VPWR VPWR hold156/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold167 hold167/A VGND VGND VPWR VPWR hold167/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold178 hold178/A VGND VGND VPWR VPWR hold178/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09913_ _13482_/Q _13671_/Q _09913_/S VGND VGND VPWR VPWR _09914_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold189 hold189/A VGND VGND VPWR VPWR hold189/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_98_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09844_ _09844_/A VGND VGND VPWR VPWR _13682_/D sky130_fd_sc_hd__clkbuf_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _09775_/A VGND VGND VPWR VPWR _13675_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06987_ _06996_/A _06996_/B VGND VGND VPWR VPWR _06987_/Y sky130_fd_sc_hd__nor2_1
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ _08728_/A _08741_/B VGND VGND VPWR VPWR _08726_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05938_ _11429_/A VGND VGND VPWR VPWR _11382_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ _08657_/A _08657_/B VGND VGND VPWR VPWR _08657_/X sky130_fd_sc_hd__or2_1
XFILLER_14_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _07645_/A _07721_/A _07627_/C VGND VGND VPWR VPWR _07610_/A sky130_fd_sc_hd__and3_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08588_ _08590_/A _08590_/B _08622_/B VGND VGND VPWR VPWR _08589_/B sky130_fd_sc_hd__a21o_1
XFILLER_41_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07539_ _07537_/Y _07538_/X _07475_/X VGND VGND VPWR VPWR _13155_/D sky130_fd_sc_hd__a21o_1
XFILLER_22_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10550_ _10562_/A _10550_/B VGND VGND VPWR VPWR _10553_/A sky130_fd_sc_hd__or2_1
X_09209_ _09210_/A _09210_/B _09220_/C VGND VGND VPWR VPWR _09214_/B sky130_fd_sc_hd__a21o_1
X_10481_ _10481_/A _10481_/B VGND VGND VPWR VPWR _10490_/B sky130_fd_sc_hd__nor2_1
X_12220_ _14124_/Q _14125_/Q _12220_/C VGND VGND VPWR VPWR _12220_/X sky130_fd_sc_hd__and3_1
XFILLER_136_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12151_ _12185_/A VGND VGND VPWR VPWR _12202_/S sky130_fd_sc_hd__buf_2
XFILLER_118_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11102_ _11065_/X _11099_/X _11101_/X _11086_/X VGND VGND VPWR VPWR _11102_/X sky130_fd_sc_hd__o211a_1
XFILLER_123_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12082_ _12082_/A VGND VGND VPWR VPWR _14458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11033_ _11033_/A VGND VGND VPWR VPWR _11033_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12984_ _13574_/CLK hold284/X VGND VGND VPWR VPWR _12984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14723_ _14724_/CLK _14723_/D VGND VGND VPWR VPWR _14723_/Q sky130_fd_sc_hd__dfxtp_1
X_11935_ _11935_/A VGND VGND VPWR VPWR _14273_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ _14709_/CLK _14654_/D VGND VGND VPWR VPWR _14654_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _11877_/A VGND VGND VPWR VPWR _11875_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _13605_/CLK _13605_/D repeater57/X VGND VGND VPWR VPWR _13605_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_60_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10817_ _10817_/A VGND VGND VPWR VPWR _13070_/D sky130_fd_sc_hd__clkbuf_1
X_14585_ _14688_/CLK _14585_/D VGND VGND VPWR VPWR hold216/A sky130_fd_sc_hd__dfxtp_1
X_11797_ _11819_/A VGND VGND VPWR VPWR _11806_/B sky130_fd_sc_hd__clkbuf_1
X_13536_ _13558_/CLK _13536_/D _12609_/A VGND VGND VPWR VPWR _13536_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10748_ _12908_/Q _10748_/B VGND VGND VPWR VPWR _10749_/A sky130_fd_sc_hd__and2_1
XFILLER_118_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13467_ _13621_/CLK _13467_/D repeater56/X VGND VGND VPWR VPWR _13467_/Q sky130_fd_sc_hd__dfrtp_1
X_10679_ _10679_/A _10687_/B VGND VGND VPWR VPWR _10680_/A sky130_fd_sc_hd__and2_1
X_12418_ _12418_/A _12418_/B input4/X VGND VGND VPWR VPWR _12419_/A sky130_fd_sc_hd__and3_1
X_13398_ _13596_/CLK hold415/X VGND VGND VPWR VPWR _13398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12349_ _14598_/Q _11959_/X _12353_/S VGND VGND VPWR VPWR _12350_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14019_ _14539_/CLK _14019_/D VGND VGND VPWR VPWR _14019_/Q sky130_fd_sc_hd__dfxtp_1
X_06910_ _13016_/Q _07968_/B VGND VGND VPWR VPWR _06919_/A sky130_fd_sc_hd__nand2_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07890_ _07898_/A _07890_/B VGND VGND VPWR VPWR _07893_/A sky130_fd_sc_hd__nand2_1
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06841_ _06852_/A _06841_/B VGND VGND VPWR VPWR _06841_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09560_ _13613_/Q _13614_/Q _13615_/Q _13616_/Q _09563_/B VGND VGND VPWR VPWR _09560_/X
+ sky130_fd_sc_hd__o41a_1
X_06772_ _07853_/B _07853_/C VGND VGND VPWR VPWR _06773_/A sky130_fd_sc_hd__and2_1
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08511_ _08481_/A _08477_/Y _08480_/B _08497_/Y VGND VGND VPWR VPWR _08512_/C sky130_fd_sc_hd__o211a_1
XFILLER_82_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09491_ _09500_/A _09491_/B VGND VGND VPWR VPWR _09509_/B sky130_fd_sc_hd__nand2_1
XFILLER_36_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08442_ _08442_/A VGND VGND VPWR VPWR _08535_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08373_ _13084_/Q _13365_/Q _08373_/S VGND VGND VPWR VPWR _08374_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07324_ _07324_/A VGND VGND VPWR VPWR _13136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07255_ _07255_/A _07255_/B VGND VGND VPWR VPWR _07258_/A sky130_fd_sc_hd__or2_1
XFILLER_137_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06206_ _14423_/Q _14421_/Q _10194_/A VGND VGND VPWR VPWR _06206_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07186_ _07186_/A VGND VGND VPWR VPWR _13349_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06137_ _06136_/X _06133_/X _10106_/A VGND VGND VPWR VPWR _06138_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06068_ _06068_/A VGND VGND VPWR VPWR _13921_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_2_0_clk clkbuf_2_3_0_clk/A VGND VGND VPWR VPWR clkbuf_3_5_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09827_ _09836_/A _09827_/B _09836_/D VGND VGND VPWR VPWR _09829_/B sky130_fd_sc_hd__and3_1
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09758_ _09758_/A _09758_/B _09758_/C VGND VGND VPWR VPWR _09760_/B sky130_fd_sc_hd__and3_1
XFILLER_74_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08709_ _08709_/A _08709_/B _08714_/D VGND VGND VPWR VPWR _08709_/Y sky130_fd_sc_hd__nand3_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _13710_/Q VGND VGND VPWR VPWR _09787_/S sky130_fd_sc_hd__inv_2
XFILLER_15_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _11720_/A VGND VGND VPWR VPWR _14052_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _14001_/Q _11519_/X _11653_/S VGND VGND VPWR VPWR _11652_/A sky130_fd_sc_hd__mux2_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10602_ _10602_/A VGND VGND VPWR VPWR _13818_/D sky130_fd_sc_hd__clkbuf_1
X_14370_ _14425_/CLK _14370_/D VGND VGND VPWR VPWR _14370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11582_ _11582_/A VGND VGND VPWR VPWR _13872_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13321_ _14742_/CLK _13321_/D VGND VGND VPWR VPWR _13321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10533_ _10533_/A _10533_/B VGND VGND VPWR VPWR _10533_/X sky130_fd_sc_hd__xor2_1
XFILLER_13_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13252_ _14690_/CLK _13252_/D hold1/X VGND VGND VPWR VPWR _13252_/Q sky130_fd_sc_hd__dfrtp_1
X_10464_ _10465_/A _10465_/B VGND VGND VPWR VPWR _10466_/A sky130_fd_sc_hd__and2_1
X_12203_ _12203_/A VGND VGND VPWR VPWR _14512_/D sky130_fd_sc_hd__clkbuf_1
X_13183_ _13423_/CLK _13183_/D VGND VGND VPWR VPWR hold367/A sky130_fd_sc_hd__dfxtp_1
X_10395_ _10396_/A _10411_/A VGND VGND VPWR VPWR _10397_/A sky130_fd_sc_hd__and2_1
XFILLER_123_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12134_ _12134_/A VGND VGND VPWR VPWR _14481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12065_ _12076_/A VGND VGND VPWR VPWR _12074_/S sky130_fd_sc_hd__buf_2
XFILLER_49_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11016_ _10991_/X _11009_/X _11014_/X _11015_/X VGND VGND VPWR VPWR _11016_/X sky130_fd_sc_hd__o211a_1
XFILLER_77_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12967_ _13265_/CLK hold369/X VGND VGND VPWR VPWR _12967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14706_ _14707_/CLK _14706_/D VGND VGND VPWR VPWR _14706_/Q sky130_fd_sc_hd__dfxtp_1
X_11918_ _14266_/Q _11478_/X _11918_/S VGND VGND VPWR VPWR _11919_/A sky130_fd_sc_hd__mux2_1
X_12898_ _12974_/CLK _12898_/D hold1/X VGND VGND VPWR VPWR _12898_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11849_ _14223_/Q _11456_/X _11853_/S VGND VGND VPWR VPWR _11850_/A sky130_fd_sc_hd__mux2_1
X_14637_ _14690_/CLK hold40/X VGND VGND VPWR VPWR _14637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14568_ _14602_/CLK _14568_/D VGND VGND VPWR VPWR _14568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13519_ _13520_/CLK _13519_/D VGND VGND VPWR VPWR _13519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14499_ _14602_/CLK _14499_/D VGND VGND VPWR VPWR _14499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07040_ _07040_/A _07165_/A VGND VGND VPWR VPWR _07059_/A sky130_fd_sc_hd__nand2_1
XFILLER_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08991_ _08951_/C _08991_/B _08991_/C VGND VGND VPWR VPWR _08995_/A sky130_fd_sc_hd__and3b_1
XFILLER_87_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07942_ _13271_/Q _07968_/B VGND VGND VPWR VPWR _07949_/D sky130_fd_sc_hd__xnor2_1
X_07873_ _07892_/A _07892_/B _07892_/C VGND VGND VPWR VPWR _07881_/B sky130_fd_sc_hd__or3_1
XFILLER_110_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09612_ _13403_/Q _13601_/Q _09620_/S VGND VGND VPWR VPWR _09613_/A sky130_fd_sc_hd__mux2_2
XFILLER_68_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06824_ _06825_/C _06823_/X VGND VGND VPWR VPWR _06824_/X sky130_fd_sc_hd__or2b_1
XFILLER_55_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09543_ _13613_/Q _09581_/B _09548_/A _09547_/A VGND VGND VPWR VPWR _09544_/B sky130_fd_sc_hd__a22o_1
XFILLER_83_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06755_ _06770_/A _06753_/A _06753_/B _06753_/C VGND VGND VPWR VPWR _07846_/C sky130_fd_sc_hd__a31o_1
XFILLER_36_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09474_ _09475_/A _09475_/B _09477_/B VGND VGND VPWR VPWR _09474_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06686_ _06665_/X _06681_/X _06682_/Y _06685_/X VGND VGND VPWR VPWR _13000_/D sky130_fd_sc_hd__a31o_1
XFILLER_24_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08425_ _08997_/A VGND VGND VPWR VPWR _13473_/D sky130_fd_sc_hd__clkbuf_2
X_08356_ _13076_/Q _13357_/Q _08362_/S VGND VGND VPWR VPWR _08357_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07307_ _07455_/A _09113_/B VGND VGND VPWR VPWR _07307_/X sky130_fd_sc_hd__and2_1
X_08287_ _08287_/A VGND VGND VPWR VPWR _13369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07238_ _08303_/A VGND VGND VPWR VPWR _08296_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_146_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07169_ _07205_/A _07205_/B VGND VGND VPWR VPWR _07174_/A sky130_fd_sc_hd__xnor2_1
XFILLER_117_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10180_ _10176_/X _10179_/X _10182_/S VGND VGND VPWR VPWR _10181_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13870_ _14656_/CLK _13870_/D VGND VGND VPWR VPWR _13870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12821_ _13653_/CLK _12821_/D VGND VGND VPWR VPWR hold161/A sky130_fd_sc_hd__dfxtp_1
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ _13702_/CLK _12752_/D VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__dfxtp_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _11703_/A VGND VGND VPWR VPWR _14033_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _13296_/CLK _12683_/D VGND VGND VPWR VPWR hold307/A sky130_fd_sc_hd__dfxtp_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _14424_/CLK _14422_/D VGND VGND VPWR VPWR _14422_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11634_ _13993_/Q _11494_/X _11634_/S VGND VGND VPWR VPWR _11635_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14353_ _14357_/CLK _14353_/D VGND VGND VPWR VPWR hold227/A sky130_fd_sc_hd__dfxtp_1
X_11565_ _11576_/A VGND VGND VPWR VPWR _11574_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_128_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13304_ _13304_/CLK hold189/X VGND VGND VPWR VPWR _13304_/Q sky130_fd_sc_hd__dfxtp_1
X_10516_ _12991_/D VGND VGND VPWR VPWR _10555_/B sky130_fd_sc_hd__inv_2
X_14284_ _14294_/CLK _14284_/D VGND VGND VPWR VPWR _14284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11496_ _11496_/A VGND VGND VPWR VPWR _13833_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13235_ _13606_/CLK hold66/X VGND VGND VPWR VPWR _13235_/Q sky130_fd_sc_hd__dfxtp_1
X_10447_ _10441_/A _10495_/A _10438_/B _10483_/B VGND VGND VPWR VPWR _10450_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_124_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13166_ _13535_/CLK _13166_/D VGND VGND VPWR VPWR hold487/A sky130_fd_sc_hd__dfxtp_1
X_10378_ _10378_/A _10378_/B VGND VGND VPWR VPWR _10378_/X sky130_fd_sc_hd__and2_1
X_12117_ _14474_/Q _11981_/X _12117_/S VGND VGND VPWR VPWR _12118_/A sky130_fd_sc_hd__mux2_1
X_13097_ _14555_/CLK hold139/X VGND VGND VPWR VPWR _13097_/Q sky130_fd_sc_hd__dfxtp_1
X_12048_ _11288_/X _14443_/Q _12052_/S VGND VGND VPWR VPWR _12049_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13999_ _14724_/CLK _13999_/D VGND VGND VPWR VPWR _13999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06540_ _06534_/B _06538_/Y _06599_/A VGND VGND VPWR VPWR _06541_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06471_ _06471_/A _06471_/B _06471_/C VGND VGND VPWR VPWR _06473_/B sky130_fd_sc_hd__and3_1
X_08210_ _13362_/Q _08210_/B VGND VGND VPWR VPWR _08211_/B sky130_fd_sc_hd__nor2_1
X_09190_ _09190_/A _09190_/B VGND VGND VPWR VPWR _09190_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08141_ _14011_/Q _14009_/Q _08161_/S VGND VGND VPWR VPWR _08141_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08072_ _08072_/A VGND VGND VPWR VPWR _12696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07023_ _10647_/B _07020_/Y _10647_/A VGND VGND VPWR VPWR _07024_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08974_ _08974_/A VGND VGND VPWR VPWR _14252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_102_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_07925_ _07925_/A _07949_/A VGND VGND VPWR VPWR _07925_/Y sky130_fd_sc_hd__nand2_1
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07856_ _07847_/A _07856_/B _13258_/Q VGND VGND VPWR VPWR _07859_/B sky130_fd_sc_hd__and3b_1
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06807_ _06807_/A VGND VGND VPWR VPWR _07876_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07787_ _07787_/A _07787_/B _07787_/C VGND VGND VPWR VPWR _07788_/B sky130_fd_sc_hd__and3_1
XFILLER_43_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09526_ _09532_/A _09526_/B VGND VGND VPWR VPWR _09534_/C sky130_fd_sc_hd__or2_1
XFILLER_83_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06738_ _07838_/B VGND VGND VPWR VPWR _07856_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09457_ _13602_/Q _09457_/B _09457_/C VGND VGND VPWR VPWR _09467_/A sky130_fd_sc_hd__and3_1
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06669_ _13038_/Q VGND VGND VPWR VPWR _06783_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_12_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08408_ _13468_/D VGND VGND VPWR VPWR _09323_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09388_ _13592_/Q _09388_/B VGND VGND VPWR VPWR _09391_/A sky130_fd_sc_hd__nor2_1
X_08339_ _08333_/A _08340_/D _08338_/Y VGND VGND VPWR VPWR _13383_/D sky130_fd_sc_hd__a21oi_1
XFILLER_137_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11350_ _11350_/A VGND VGND VPWR VPWR _13773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10301_ _14639_/Q _14640_/Q _14646_/Q _12336_/C VGND VGND VPWR VPWR _10302_/A sky130_fd_sc_hd__or4_1
XFILLER_137_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11281_ _11330_/A VGND VGND VPWR VPWR _11376_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_118_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13020_ _13031_/CLK _13020_/D repeater59/X VGND VGND VPWR VPWR _13020_/Q sky130_fd_sc_hd__dfrtp_1
X_10232_ _14522_/D _10231_/X _14557_/D VGND VGND VPWR VPWR _10233_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10163_ _10163_/A VGND VGND VPWR VPWR _14119_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10094_ _10094_/A VGND VGND VPWR VPWR _13906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13922_ _14047_/CLK hold213/X VGND VGND VPWR VPWR _13922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13853_ _14180_/CLK _13853_/D VGND VGND VPWR VPWR _13853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12804_ _14108_/CLK _12804_/D VGND VGND VPWR VPWR hold347/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10996_ _14299_/Q _14469_/Q _14225_/Q _14055_/Q _10993_/X _10995_/X VGND VGND VPWR
+ VPWR _10996_/X sky130_fd_sc_hd__mux4_1
X_13784_ _13945_/CLK _13784_/D VGND VGND VPWR VPWR _13784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _14696_/CLK _12735_/D VGND VGND VPWR VPWR hold470/A sky130_fd_sc_hd__dfxtp_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _14678_/CLK _12666_/D VGND VGND VPWR VPWR _13247_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11617_ _13985_/Q _11469_/X _11623_/S VGND VGND VPWR VPWR _11618_/A sky130_fd_sc_hd__mux2_1
X_14405_ _14410_/CLK _14405_/D VGND VGND VPWR VPWR _14405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12597_ _10901_/X hold344/X _12580_/X VGND VGND VPWR VPWR _14729_/D sky130_fd_sc_hd__o21a_1
XFILLER_7_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11548_ _13633_/Q _11552_/B VGND VGND VPWR VPWR _11549_/A sky130_fd_sc_hd__and2_1
X_14336_ _14557_/CLK _14336_/D VGND VGND VPWR VPWR hold217/A sky130_fd_sc_hd__dfxtp_1
XFILLER_143_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold508 hold508/A VGND VGND VPWR VPWR hold508/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold519 hold519/A VGND VGND VPWR VPWR hold519/X sky130_fd_sc_hd__clkbuf_2
X_14267_ _14714_/CLK _14267_/D VGND VGND VPWR VPWR _14267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11479_ _13828_/Q _11478_/X _11479_/S VGND VGND VPWR VPWR _11480_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13218_ _13423_/CLK hold376/X VGND VGND VPWR VPWR _13218_/Q sky130_fd_sc_hd__dfxtp_1
X_14198_ _14210_/CLK _14198_/D VGND VGND VPWR VPWR _14198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13149_ _13555_/CLK _13149_/D repeater57/X VGND VGND VPWR VPWR _13149_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05971_ _13625_/Q _13626_/Q _13627_/Q _13628_/Q VGND VGND VPWR VPWR _05977_/A sky130_fd_sc_hd__or4_1
XFILLER_100_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07710_ _07733_/B _07710_/B _07710_/C VGND VGND VPWR VPWR _07735_/A sky130_fd_sc_hd__and3_1
X_08690_ _13451_/Q _09576_/B _08689_/X VGND VGND VPWR VPWR _08698_/A sky130_fd_sc_hd__a21oi_1
XFILLER_38_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07641_ _07641_/A _07641_/B _07656_/B VGND VGND VPWR VPWR _07654_/A sky130_fd_sc_hd__or3_1
XFILLER_38_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07572_ _13160_/Q _09277_/B VGND VGND VPWR VPWR _07572_/X sky130_fd_sc_hd__or2_1
XFILLER_15_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09311_ _09311_/A VGND VGND VPWR VPWR _12783_/D sky130_fd_sc_hd__clkbuf_1
X_06523_ _06563_/B _06524_/C VGND VGND VPWR VPWR _06525_/B sky130_fd_sc_hd__and2_1
XFILLER_22_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09242_ _09242_/A _09242_/B _09242_/C _09242_/D VGND VGND VPWR VPWR _09242_/X sky130_fd_sc_hd__or4_1
X_06454_ _06454_/A VGND VGND VPWR VPWR _12880_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09173_ _09173_/A _09173_/B VGND VGND VPWR VPWR _09174_/B sky130_fd_sc_hd__nand2_1
X_06385_ _06455_/A _06444_/A VGND VGND VPWR VPWR _06429_/B sky130_fd_sc_hd__and2b_1
XFILLER_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08124_ _08124_/A _08124_/B VGND VGND VPWR VPWR _08124_/X sky130_fd_sc_hd__and2_1
XFILLER_107_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08055_ _08055_/A VGND VGND VPWR VPWR _12688_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07006_ _07003_/Y _07004_/X _06999_/A _07005_/Y VGND VGND VPWR VPWR _07006_/X sky130_fd_sc_hd__a211o_1
XFILLER_162_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput39 _13336_/Q VGND VGND VPWR VPWR data_o[18] sky130_fd_sc_hd__buf_2
XFILLER_163_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08957_ _08993_/A _08993_/B VGND VGND VPWR VPWR _08962_/A sky130_fd_sc_hd__xnor2_1
XFILLER_56_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07908_ _07914_/B _07907_/Y _06859_/X VGND VGND VPWR VPWR _13266_/D sky130_fd_sc_hd__a21o_1
X_08888_ _08919_/A _08919_/B VGND VGND VPWR VPWR _08889_/B sky130_fd_sc_hd__xnor2_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07839_ _13257_/Q _07840_/B VGND VGND VPWR VPWR _07839_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10850_ _13143_/Q _10852_/B VGND VGND VPWR VPWR _10851_/A sky130_fd_sc_hd__and2_1
XFILLER_71_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09509_ _09509_/A _09509_/B _09509_/C _09509_/D VGND VGND VPWR VPWR _09535_/A sky130_fd_sc_hd__or4_1
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10781_ _10781_/A VGND VGND VPWR VPWR _10790_/B sky130_fd_sc_hd__clkbuf_1
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12520_ _12520_/A VGND VGND VPWR VPWR _14706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _12451_/A VGND VGND VPWR VPWR _14657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11402_ _11402_/A VGND VGND VPWR VPWR _13793_/D sky130_fd_sc_hd__clkbuf_1
X_12382_ _14613_/Q _12007_/X _12386_/S VGND VGND VPWR VPWR _12383_/A sky130_fd_sc_hd__mux2_1
XANTENNA_90 _13091_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14121_ _14159_/CLK hold308/X VGND VGND VPWR VPWR _14121_/Q sky130_fd_sc_hd__dfxtp_1
X_11333_ _13878_/Q _13844_/Q VGND VGND VPWR VPWR _11364_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14052_ _14704_/CLK _14052_/D VGND VGND VPWR VPWR _14052_/Q sky130_fd_sc_hd__dfxtp_1
X_11264_ _12626_/B _11264_/B VGND VGND VPWR VPWR _11264_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13003_ _13256_/CLK _13003_/D hold1/X VGND VGND VPWR VPWR _13003_/Q sky130_fd_sc_hd__dfrtp_1
X_10215_ _10215_/A VGND VGND VPWR VPWR _14395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11195_ _13335_/Q _11150_/X _11184_/X _11194_/Y VGND VGND VPWR VPWR _13335_/D sky130_fd_sc_hd__o22a_1
XFILLER_79_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10146_ _10146_/A VGND VGND VPWR VPWR _14287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10077_ _10016_/A _10057_/X _10072_/X VGND VGND VPWR VPWR _10077_/X sky130_fd_sc_hd__a21o_1
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13905_ _14693_/CLK _13905_/D VGND VGND VPWR VPWR hold331/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13836_ _14721_/CLK _13836_/D VGND VGND VPWR VPWR _13836_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10979_ _13320_/Q _10907_/X _10967_/X _10978_/Y VGND VGND VPWR VPWR _13320_/D sky130_fd_sc_hd__o22a_1
X_13767_ _14717_/CLK _13767_/D VGND VGND VPWR VPWR _13767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12718_ _13366_/CLK _12718_/D VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__dfxtp_1
XFILLER_149_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13698_ _13698_/CLK _13698_/D repeater57/X VGND VGND VPWR VPWR _13698_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_129_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12649_ _14749_/Q _12649_/B VGND VGND VPWR VPWR _12649_/X sky130_fd_sc_hd__or2_1
XFILLER_129_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06170_ _06170_/A VGND VGND VPWR VPWR _14172_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14319_ _14319_/CLK hold173/X VGND VGND VPWR VPWR hold77/A sky130_fd_sc_hd__dfxtp_2
Xhold305 hold305/A VGND VGND VPWR VPWR hold305/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold316 hold316/A VGND VGND VPWR VPWR hold316/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold327 hold327/A VGND VGND VPWR VPWR hold327/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold338 hold338/A VGND VGND VPWR VPWR hold338/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold349 hold349/A VGND VGND VPWR VPWR hold349/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09860_ _13685_/Q _09851_/A _09858_/D _13686_/Q VGND VGND VPWR VPWR _09861_/C sky130_fd_sc_hd__a31o_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _11268_/B _08808_/Y _11268_/A VGND VGND VPWR VPWR _08812_/A sky130_fd_sc_hd__mux2_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09791_ _13677_/Q _09791_/B VGND VGND VPWR VPWR _09804_/A sky130_fd_sc_hd__nor2_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08742_ _08742_/A _08742_/B VGND VGND VPWR VPWR _08742_/Y sky130_fd_sc_hd__nor2_1
X_05954_ _06309_/S VGND VGND VPWR VPWR _06313_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08673_ _09518_/B VGND VGND VPWR VPWR _08730_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_26_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_186_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _14619_/CLK sky130_fd_sc_hd__clkbuf_16
X_07624_ _07723_/B VGND VGND VPWR VPWR _07745_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07555_ _13158_/Q _09270_/B VGND VGND VPWR VPWR _07559_/B sky130_fd_sc_hd__xnor2_1
XFILLER_81_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06506_ _06506_/A _06516_/A VGND VGND VPWR VPWR _06508_/A sky130_fd_sc_hd__or2_1
XFILLER_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07486_ _07499_/A VGND VGND VPWR VPWR _07486_/X sky130_fd_sc_hd__buf_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09225_ _09226_/B _09224_/X _07526_/X VGND VGND VPWR VPWR _13543_/D sky130_fd_sc_hd__o21bai_1
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06437_ _06437_/A _06437_/B VGND VGND VPWR VPWR _06437_/X sky130_fd_sc_hd__xor2_1
XFILLER_148_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09156_ _09156_/A _09156_/B _09156_/C VGND VGND VPWR VPWR _09156_/Y sky130_fd_sc_hd__nand3_1
X_06368_ _06368_/A VGND VGND VPWR VPWR _13754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08107_ _13424_/Q VGND VGND VPWR VPWR _08142_/A sky130_fd_sc_hd__clkbuf_2
X_09087_ _07261_/B _09086_/C _13524_/Q VGND VGND VPWR VPWR _09089_/B sky130_fd_sc_hd__a21oi_1
X_06299_ _13870_/Q _13854_/Q _06309_/S VGND VGND VPWR VPWR _06300_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_110_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _13610_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_163_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08038_ _12957_/Q _13257_/Q _08040_/S VGND VGND VPWR VPWR _08039_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10000_ _10000_/A VGND VGND VPWR VPWR _12667_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09989_ _09989_/A VGND VGND VPWR VPWR _13707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11951_ _12342_/A _12095_/B VGND VGND VPWR VPWR _12001_/A sky130_fd_sc_hd__nor2_4
Xclkbuf_leaf_177_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _14652_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10902_ input28/X VGND VGND VPWR VPWR _12596_/B sky130_fd_sc_hd__inv_2
X_11882_ _14238_/Q _11504_/X _11886_/S VGND VGND VPWR VPWR _11883_/A sky130_fd_sc_hd__mux2_1
X_14670_ _14704_/CLK _14670_/D VGND VGND VPWR VPWR _14670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13621_ _13621_/CLK _13621_/D repeater56/X VGND VGND VPWR VPWR _13621_/Q sky130_fd_sc_hd__dfrtp_1
X_10833_ _13135_/Q _10841_/B VGND VGND VPWR VPWR _10834_/A sky130_fd_sc_hd__and2_1
XFILLER_72_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13552_ _13552_/CLK _13552_/D _12609_/A VGND VGND VPWR VPWR _13552_/Q sky130_fd_sc_hd__dfrtp_4
X_10764_ _13004_/Q _10768_/B VGND VGND VPWR VPWR _10765_/A sky130_fd_sc_hd__and2_1
XFILLER_13_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater58 hold1/X VGND VGND VPWR VPWR _12609_/A sky130_fd_sc_hd__buf_12
X_12503_ _12503_/A VGND VGND VPWR VPWR _14689_/D sky130_fd_sc_hd__clkbuf_1
X_13483_ _14251_/CLK hold195/X VGND VGND VPWR VPWR _13483_/Q sky130_fd_sc_hd__dfxtp_1
X_10695_ _10695_/A VGND VGND VPWR VPWR _12926_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12434_ _12434_/A VGND VGND VPWR VPWR _14649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12365_ _12365_/A VGND VGND VPWR VPWR _14605_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_101_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _13805_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11316_ _11316_/A VGND VGND VPWR VPWR _13765_/D sky130_fd_sc_hd__clkbuf_1
X_14104_ _14410_/CLK _14104_/D VGND VGND VPWR VPWR _14104_/Q sky130_fd_sc_hd__dfxtp_1
X_12296_ _14564_/Q _11972_/X _12302_/S VGND VGND VPWR VPWR _12297_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14035_ _14725_/CLK _14035_/D VGND VGND VPWR VPWR _14035_/Q sky130_fd_sc_hd__dfxtp_1
X_11247_ _11207_/X _11244_/X _11246_/X _12647_/A VGND VGND VPWR VPWR _11247_/X sky130_fd_sc_hd__o211a_1
XFILLER_106_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11178_ _11159_/X _11175_/Y _11177_/Y _11166_/X VGND VGND VPWR VPWR _11179_/B sky130_fd_sc_hd__a211o_1
X_10129_ _13865_/Q _13849_/Q _14167_/D VGND VGND VPWR VPWR _10130_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_168_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _14425_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_82_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13819_ _14533_/CLK _13819_/D VGND VGND VPWR VPWR _13819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07340_ _07318_/B _07322_/B _07337_/Y _07316_/A VGND VGND VPWR VPWR _07341_/B sky130_fd_sc_hd__o211a_1
XFILLER_32_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07271_ _07231_/Y _07388_/B _07270_/X _07228_/X VGND VGND VPWR VPWR _07284_/B sky130_fd_sc_hd__a22oi_4
XFILLER_148_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09010_ _13206_/Q _13435_/Q _09018_/S VGND VGND VPWR VPWR _09011_/A sky130_fd_sc_hd__mux2_1
X_06222_ _14399_/Q _14391_/Q _06321_/S VGND VGND VPWR VPWR _06222_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06153_ _10616_/A _06152_/X _10121_/S VGND VGND VPWR VPWR _06154_/A sky130_fd_sc_hd__mux2_1
Xhold102 hold102/A VGND VGND VPWR VPWR hold102/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_117_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold113 hold113/A VGND VGND VPWR VPWR hold113/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_145_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold124 hold124/A VGND VGND VPWR VPWR hold124/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold135 hold135/A VGND VGND VPWR VPWR hold135/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_117_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06084_ _06084_/A VGND VGND VPWR VPWR _13966_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold146 hold146/A VGND VGND VPWR VPWR hold146/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold157 hold157/A VGND VGND VPWR VPWR hold157/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold168 hold168/A VGND VGND VPWR VPWR hold168/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09912_ _09912_/A VGND VGND VPWR VPWR _12844_/D sky130_fd_sc_hd__clkbuf_1
Xhold179 hold179/A VGND VGND VPWR VPWR hold179/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09843_ _09838_/B _09842_/Y _09855_/A VGND VGND VPWR VPWR _09844_/A sky130_fd_sc_hd__mux2_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06986_ _06986_/A _06986_/B VGND VGND VPWR VPWR _06996_/B sky130_fd_sc_hd__or2_1
XFILLER_86_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09774_ _09769_/B _09773_/Y _09774_/S VGND VGND VPWR VPWR _09775_/A sky130_fd_sc_hd__mux2_1
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08725_ _08728_/A _08741_/B VGND VGND VPWR VPWR _08725_/X sky130_fd_sc_hd__or2_1
X_05937_ _05937_/A _05937_/B VGND VGND VPWR VPWR _11429_/A sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_159_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _14710_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _08617_/X _08652_/Y _08664_/B _08655_/X VGND VGND VPWR VPWR _13449_/D sky130_fd_sc_hd__a31o_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07607_ _13245_/D VGND VGND VPWR VPWR _07721_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _08587_/A _08621_/A VGND VGND VPWR VPWR _08622_/B sky130_fd_sc_hd__or2_1
X_07538_ _07548_/A _07547_/A _08296_/B VGND VGND VPWR VPWR _07538_/X sky130_fd_sc_hd__o21a_1
X_07469_ _09258_/B VGND VGND VPWR VPWR _09270_/B sky130_fd_sc_hd__clkbuf_2
X_09208_ _09214_/A _09208_/B VGND VGND VPWR VPWR _09220_/C sky130_fd_sc_hd__nand2_1
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10480_ _10480_/A _10480_/B VGND VGND VPWR VPWR _10490_/A sky130_fd_sc_hd__nor2_1
XFILLER_108_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09139_ _13532_/Q _09139_/B _09139_/C VGND VGND VPWR VPWR _09161_/B sky130_fd_sc_hd__and3_1
XFILLER_136_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12150_ _12150_/A _12342_/B VGND VGND VPWR VPWR _12185_/A sky130_fd_sc_hd__nor2_4
XFILLER_136_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11101_ _11101_/A _11084_/X VGND VGND VPWR VPWR _11101_/X sky130_fd_sc_hd__or2b_1
XFILLER_151_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12081_ _11343_/X _14458_/Q _12085_/S VGND VGND VPWR VPWR _12082_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11032_ _14602_/Q _14564_/Q _14495_/Q _14447_/Q _10969_/X _10970_/X VGND VGND VPWR
+ VPWR _11033_/A sky130_fd_sc_hd__mux4_1
XFILLER_1_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12983_ _13274_/CLK hold333/X VGND VGND VPWR VPWR _12983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14722_ _14722_/CLK _14722_/D VGND VGND VPWR VPWR _14722_/Q sky130_fd_sc_hd__dfxtp_1
X_11934_ _14273_/Q _11501_/X _11940_/S VGND VGND VPWR VPWR _11935_/A sky130_fd_sc_hd__mux2_1
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14653_ _14710_/CLK _14653_/D VGND VGND VPWR VPWR _14653_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _11865_/A VGND VGND VPWR VPWR _14230_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13604_ _13604_/CLK _13604_/D repeater56/X VGND VGND VPWR VPWR _13604_/Q sky130_fd_sc_hd__dfrtp_1
X_10816_ _13028_/Q _10818_/B VGND VGND VPWR VPWR _10817_/A sky130_fd_sc_hd__and2_1
X_14584_ _14688_/CLK hold216/X VGND VGND VPWR VPWR _14584_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_158_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11796_ _11796_/A VGND VGND VPWR VPWR _14091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13535_ _13535_/CLK _13535_/D repeater57/X VGND VGND VPWR VPWR _13535_/Q sky130_fd_sc_hd__dfrtp_1
X_10747_ _10747_/A VGND VGND VPWR VPWR _12950_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13466_ _13622_/CLK _13466_/D repeater57/X VGND VGND VPWR VPWR _13466_/Q sky130_fd_sc_hd__dfrtp_1
X_10678_ _10748_/B VGND VGND VPWR VPWR _10687_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_145_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12417_ _12417_/A VGND VGND VPWR VPWR _14642_/D sky130_fd_sc_hd__clkbuf_1
X_13397_ _13596_/CLK hold483/X VGND VGND VPWR VPWR _13397_/Q sky130_fd_sc_hd__dfxtp_1
X_12348_ _12348_/A VGND VGND VPWR VPWR _14597_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12279_ _12279_/A VGND VGND VPWR VPWR _14554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14018_ _14357_/CLK _14018_/D VGND VGND VPWR VPWR _14018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06840_ _06840_/A VGND VGND VPWR VPWR _07895_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_56_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06771_ _06719_/A _06786_/B _06770_/C VGND VGND VPWR VPWR _07853_/C sky130_fd_sc_hd__a21o_1
XFILLER_83_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08510_ _13439_/Q _09394_/B VGND VGND VPWR VPWR _08512_/B sky130_fd_sc_hd__xnor2_1
X_09490_ _13606_/Q _09518_/B VGND VGND VPWR VPWR _09491_/B sky130_fd_sc_hd__or2_1
XFILLER_63_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08441_ _13471_/Q VGND VGND VPWR VPWR _08442_/A sky130_fd_sc_hd__inv_2
XFILLER_51_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08372_ _08372_/A VGND VGND VPWR VPWR _12719_/D sky130_fd_sc_hd__clkbuf_1
X_07323_ _09120_/B _07322_/X _09182_/A VGND VGND VPWR VPWR _07324_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07254_ _07261_/B _09086_/C _13132_/Q VGND VGND VPWR VPWR _07255_/B sky130_fd_sc_hd__a21oi_1
XFILLER_164_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06205_ _06205_/A VGND VGND VPWR VPWR _14369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07185_ _07156_/Y _07184_/X _07199_/S VGND VGND VPWR VPWR _07186_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06136_ _14206_/Q _14204_/Q _10107_/A VGND VGND VPWR VPWR _06136_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06067_ _06066_/X _06063_/X _10019_/A VGND VGND VPWR VPWR _06068_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09826_ _09826_/A VGND VGND VPWR VPWR _13680_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09757_ _09735_/A _09836_/B _14440_/Q _09778_/A VGND VGND VPWR VPWR _09758_/C sky130_fd_sc_hd__a31o_1
X_06969_ _13024_/Q _07988_/B VGND VGND VPWR VPWR _06978_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08708_ _08709_/A _08709_/B _08714_/D VGND VGND VPWR VPWR _08708_/X sky130_fd_sc_hd__a21o_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _14214_/Q _14212_/Q _09688_/S VGND VGND VPWR VPWR _09688_/X sky130_fd_sc_hd__mux2_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _08644_/A _08653_/A VGND VGND VPWR VPWR _08641_/A sky130_fd_sc_hd__or2_1
XFILLER_15_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11650_ _11650_/A VGND VGND VPWR VPWR _14000_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10601_ _10601_/A _14635_/D _10601_/C VGND VGND VPWR VPWR _10602_/A sky130_fd_sc_hd__and3_1
XFILLER_11_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11581_ _13648_/Q _11585_/B VGND VGND VPWR VPWR _11582_/A sky130_fd_sc_hd__and2_1
XFILLER_22_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10532_ _10531_/B _10532_/B VGND VGND VPWR VPWR _10533_/B sky130_fd_sc_hd__and2b_1
X_13320_ _14742_/CLK _13320_/D VGND VGND VPWR VPWR _13320_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10463_ _10463_/A _10463_/B VGND VGND VPWR VPWR _10465_/B sky130_fd_sc_hd__xor2_1
XFILLER_89_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13251_ _13596_/CLK hold99/X VGND VGND VPWR VPWR _13522_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_108_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12202_ _14512_/Q _12025_/X _12202_/S VGND VGND VPWR VPWR _12203_/A sky130_fd_sc_hd__mux2_1
X_13182_ _13423_/CLK _13182_/D VGND VGND VPWR VPWR hold493/A sky130_fd_sc_hd__dfxtp_1
X_10394_ _10407_/B _10394_/B VGND VGND VPWR VPWR _10411_/A sky130_fd_sc_hd__nor2_1
XFILLER_151_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12133_ _14481_/Q _12004_/X _12139_/S VGND VGND VPWR VPWR _12134_/A sky130_fd_sc_hd__mux2_1
X_12064_ _12064_/A VGND VGND VPWR VPWR _14450_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11015_ _11224_/A VGND VGND VPWR VPWR _11015_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12966_ _13265_/CLK hold196/X VGND VGND VPWR VPWR _12966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14705_ _14705_/CLK _14705_/D VGND VGND VPWR VPWR _14705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11917_ _11917_/A VGND VGND VPWR VPWR _14265_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _13273_/CLK _12897_/D repeater59/X VGND VGND VPWR VPWR _12897_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _14636_/CLK hold322/X VGND VGND VPWR VPWR hold123/A sky130_fd_sc_hd__dfxtp_1
X_11848_ _11848_/A VGND VGND VPWR VPWR _14222_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14567_ _14712_/CLK _14567_/D VGND VGND VPWR VPWR _14567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11779_ _11779_/A VGND VGND VPWR VPWR _14083_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13518_ _13520_/CLK _13518_/D VGND VGND VPWR VPWR _13518_/Q sky130_fd_sc_hd__dfxtp_1
X_14498_ _14712_/CLK _14498_/D VGND VGND VPWR VPWR _14498_/Q sky130_fd_sc_hd__dfxtp_1
X_13449_ _13704_/CLK _13449_/D repeater56/X VGND VGND VPWR VPWR _13449_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08990_ _08966_/A _08993_/C _08985_/A VGND VGND VPWR VPWR _08996_/A sky130_fd_sc_hd__a21o_1
X_07941_ _07909_/X _07944_/B _07939_/Y _07940_/X VGND VGND VPWR VPWR _13270_/D sky130_fd_sc_hd__a31o_1
XFILLER_96_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07872_ _07860_/A _07860_/B _07884_/C VGND VGND VPWR VPWR _07892_/C sky130_fd_sc_hd__o21a_1
XFILLER_56_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09611_ _09644_/A VGND VGND VPWR VPWR _09620_/S sky130_fd_sc_hd__clkbuf_2
X_06823_ _13008_/Q _07876_/B _06825_/B VGND VGND VPWR VPWR _06823_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09542_ _13614_/Q _09542_/B VGND VGND VPWR VPWR _09547_/B sky130_fd_sc_hd__xor2_1
X_06754_ _06770_/A _06786_/B VGND VGND VPWR VPWR _07846_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09473_ _09473_/A _09473_/B VGND VGND VPWR VPWR _09477_/B sky130_fd_sc_hd__or2_1
X_06685_ _06859_/A _07821_/B VGND VGND VPWR VPWR _06685_/X sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_90_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _13673_/CLK sky130_fd_sc_hd__clkbuf_16
X_08424_ _09002_/A VGND VGND VPWR VPWR _08997_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08355_ _08355_/A VGND VGND VPWR VPWR _12711_/D sky130_fd_sc_hd__clkbuf_1
X_07306_ _07305_/A _07305_/C _07305_/B VGND VGND VPWR VPWR _07306_/Y sky130_fd_sc_hd__o21ai_1
X_08286_ _08281_/B _08285_/Y _08286_/S VGND VGND VPWR VPWR _08287_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07237_ _09088_/B _07237_/B VGND VGND VPWR VPWR _13131_/D sky130_fd_sc_hd__xnor2_1
XFILLER_118_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07168_ _07168_/A VGND VGND VPWR VPWR _07205_/B sky130_fd_sc_hd__inv_2
XFILLER_117_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06119_ _14161_/Q _06119_/B VGND VGND VPWR VPWR _06127_/A sky130_fd_sc_hd__xnor2_2
XFILLER_105_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07099_ _07075_/A _07075_/B _07073_/B VGND VGND VPWR VPWR _07131_/B sky130_fd_sc_hd__a21oi_1
XFILLER_132_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09809_ _09836_/A _09809_/B _09809_/C VGND VGND VPWR VPWR _09811_/B sky130_fd_sc_hd__and3_1
XFILLER_46_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12820_ _13855_/CLK _12820_/D VGND VGND VPWR VPWR hold188/A sky130_fd_sc_hd__dfxtp_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12751_ _13702_/CLK _12751_/D VGND VGND VPWR VPWR hold176/A sky130_fd_sc_hd__dfxtp_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_81_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _14678_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11702_ _14033_/Q _11513_/X _11708_/S VGND VGND VPWR VPWR _11703_/A sky130_fd_sc_hd__mux2_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _13296_/CLK _12682_/D VGND VGND VPWR VPWR hold352/A sky130_fd_sc_hd__dfxtp_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14421_ _14424_/CLK _14421_/D VGND VGND VPWR VPWR _14421_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _11633_/A VGND VGND VPWR VPWR _13992_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14352_ _14357_/CLK _14352_/D VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__dfxtp_1
X_11564_ _11564_/A VGND VGND VPWR VPWR _13864_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13303_ _13303_/CLK hold105/X VGND VGND VPWR VPWR _13303_/Q sky130_fd_sc_hd__dfxtp_1
X_10515_ _12992_/D VGND VGND VPWR VPWR _10567_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14283_ _14294_/CLK _14283_/D VGND VGND VPWR VPWR _14283_/Q sky130_fd_sc_hd__dfxtp_1
X_11495_ _13833_/Q _11494_/X _11495_/S VGND VGND VPWR VPWR _11496_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10446_ _10460_/A VGND VGND VPWR VPWR _10483_/B sky130_fd_sc_hd__inv_2
X_13234_ _13617_/CLK hold426/X VGND VGND VPWR VPWR _13234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10377_ _10377_/A _10396_/A VGND VGND VPWR VPWR _10398_/B sky130_fd_sc_hd__nor2_1
XFILLER_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13165_ _13423_/CLK _13165_/D VGND VGND VPWR VPWR _13165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12116_ _12116_/A VGND VGND VPWR VPWR _14473_/D sky130_fd_sc_hd__clkbuf_1
X_13096_ _13587_/CLK hold410/X VGND VGND VPWR VPWR _13096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12047_ _12047_/A VGND VGND VPWR VPWR _14442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13998_ _14722_/CLK _13998_/D VGND VGND VPWR VPWR _13998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12949_ _13274_/CLK _12949_/D VGND VGND VPWR VPWR hold260/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_72_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _13366_/CLK sky130_fd_sc_hd__clkbuf_16
X_06470_ _06543_/A _14439_/Q _10339_/A _06482_/A VGND VGND VPWR VPWR _06471_/C sky130_fd_sc_hd__a31o_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_1_0_clk clkbuf_2_1_0_clk/A VGND VGND VPWR VPWR clkbuf_3_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_14619_ _14619_/CLK _14619_/D VGND VGND VPWR VPWR _14619_/Q sky130_fd_sc_hd__dfxtp_1
X_08140_ _08140_/A VGND VGND VPWR VPWR _13356_/D sky130_fd_sc_hd__clkbuf_1
X_08071_ _12972_/Q _13272_/Q _08073_/S VGND VGND VPWR VPWR _08072_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07022_ _07218_/S VGND VGND VPWR VPWR _10647_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08973_ _08944_/Y _08972_/X _08987_/S VGND VGND VPWR VPWR _08974_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_07924_ _07925_/A _07949_/A VGND VGND VPWR VPWR _07924_/X sky130_fd_sc_hd__or2_1
XFILLER_130_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_56_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07855_ _07885_/A _07885_/B VGND VGND VPWR VPWR _07860_/A sky130_fd_sc_hd__or2_1
X_06806_ _06825_/A _06806_/B VGND VGND VPWR VPWR _06806_/Y sky130_fd_sc_hd__nand2_1
X_07786_ _07786_/A _07786_/B VGND VGND VPWR VPWR _07788_/A sky130_fd_sc_hd__and2_1
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09525_ _13611_/Q _09525_/B VGND VGND VPWR VPWR _09526_/B sky130_fd_sc_hd__nor2_1
X_06737_ _06737_/A _06753_/B VGND VGND VPWR VPWR _07838_/B sky130_fd_sc_hd__xnor2_4
XFILLER_25_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_63_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _13256_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09456_ _09437_/X _09460_/B _09455_/Y _08631_/X VGND VGND VPWR VPWR _13601_/D sky130_fd_sc_hd__a31o_1
X_06668_ _13350_/Q _13348_/Q _06705_/S VGND VGND VPWR VPWR _06668_/X sky130_fd_sc_hd__mux2_1
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08407_ _08407_/A VGND VGND VPWR VPWR _12735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06599_ _06599_/A VGND VGND VPWR VPWR _06599_/X sky130_fd_sc_hd__clkbuf_2
X_09387_ _09387_/A VGND VGND VPWR VPWR _13592_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08338_ _08338_/A _08338_/B VGND VGND VPWR VPWR _08338_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08269_ _08338_/A _08267_/Y _08268_/Y VGND VGND VPWR VPWR _13367_/D sky130_fd_sc_hd__a21oi_1
XFILLER_137_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10300_ _14687_/Q _14688_/Q VGND VGND VPWR VPWR _14583_/D sky130_fd_sc_hd__xnor2_1
X_11280_ _12150_/A _12510_/A VGND VGND VPWR VPWR _11330_/A sky130_fd_sc_hd__nor2_8
XFILLER_125_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10231_ _14369_/Q _10230_/X _10234_/A VGND VGND VPWR VPWR _10231_/X sky130_fd_sc_hd__a21o_1
XFILLER_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10162_ _14290_/D _10161_/X _14292_/D VGND VGND VPWR VPWR _10163_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10093_ _10089_/X _10092_/X _10095_/S VGND VGND VPWR VPWR _10094_/A sky130_fd_sc_hd__mux2_1
X_13921_ _14042_/CLK _13921_/D VGND VGND VPWR VPWR _13921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13852_ _14180_/CLK _13852_/D VGND VGND VPWR VPWR _13852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12803_ _14275_/CLK _12803_/D VGND VGND VPWR VPWR hold166/A sky130_fd_sc_hd__dfxtp_1
X_13783_ _13799_/CLK _13783_/D VGND VGND VPWR VPWR _13783_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_54_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _14643_/CLK sky130_fd_sc_hd__clkbuf_16
X_10995_ _10995_/A VGND VGND VPWR VPWR _10995_/X sky130_fd_sc_hd__buf_2
XFILLER_16_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12734_ _14696_/CLK _12734_/D VGND VGND VPWR VPWR hold363/A sky130_fd_sc_hd__dfxtp_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _14678_/CLK _12665_/D VGND VGND VPWR VPWR _13246_/D sky130_fd_sc_hd__dfxtp_2
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _14410_/CLK _14404_/D VGND VGND VPWR VPWR _14404_/Q sky130_fd_sc_hd__dfxtp_1
X_11616_ _11616_/A VGND VGND VPWR VPWR _13984_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12596_ _14729_/Q _12596_/B VGND VGND VPWR VPWR hold344/A sky130_fd_sc_hd__and2_1
XFILLER_129_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14335_ _14557_/CLK hold217/X VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11547_ _11547_/A VGND VGND VPWR VPWR _13856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold509 hold509/A VGND VGND VPWR VPWR hold509/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14266_ _14657_/CLK _14266_/D VGND VGND VPWR VPWR _14266_/Q sky130_fd_sc_hd__dfxtp_1
X_11478_ _14514_/Q VGND VGND VPWR VPWR _11478_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13217_ _13621_/CLK hold518/X VGND VGND VPWR VPWR _13217_/Q sky130_fd_sc_hd__dfxtp_1
X_10429_ _10415_/C _10431_/B _10429_/C VGND VGND VPWR VPWR _10430_/A sky130_fd_sc_hd__and3b_1
XFILLER_124_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14197_ _14209_/CLK _14197_/D VGND VGND VPWR VPWR _14197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _13535_/CLK _13148_/D repeater57/X VGND VGND VPWR VPWR _13148_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05970_ _05970_/A _05970_/B _05970_/C VGND VGND VPWR VPWR _05970_/X sky130_fd_sc_hd__and3_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13079_ _13434_/CLK hold122/X VGND VGND VPWR VPWR _13079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07640_ _07633_/B _07640_/B VGND VGND VPWR VPWR _07659_/A sky130_fd_sc_hd__and2b_1
XFILLER_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07571_ _13160_/Q _07579_/B VGND VGND VPWR VPWR _07571_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_45_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _14439_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_81_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09310_ _13293_/Q _13531_/Q _09310_/S VGND VGND VPWR VPWR _09311_/A sky130_fd_sc_hd__mux2_1
X_06522_ _06522_/A VGND VGND VPWR VPWR _12886_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09241_ _09241_/A _09241_/B VGND VGND VPWR VPWR _09242_/D sky130_fd_sc_hd__nand2_1
X_06453_ _06448_/B _06452_/X _06622_/B VGND VGND VPWR VPWR _06454_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09172_ _09172_/A _09172_/B VGND VGND VPWR VPWR _09190_/A sky130_fd_sc_hd__nor2_1
X_06384_ _13108_/D VGND VGND VPWR VPWR _06444_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08123_ _08123_/A _08123_/B VGND VGND VPWR VPWR _08124_/B sky130_fd_sc_hd__xnor2_1
XFILLER_135_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08054_ _12964_/Q _13264_/Q _08062_/S VGND VGND VPWR VPWR _08055_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07005_ _07001_/B _07001_/C _07001_/A VGND VGND VPWR VPWR _07005_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_115_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08956_ _08956_/A VGND VGND VPWR VPWR _08993_/B sky130_fd_sc_hd__inv_2
XFILLER_103_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07907_ _07916_/A _07906_/B _06743_/A VGND VGND VPWR VPWR _07907_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08887_ _08863_/A _08863_/B _08861_/B VGND VGND VPWR VPWR _08919_/B sky130_fd_sc_hd__a21oi_1
XFILLER_17_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07838_ _13258_/Q _07838_/B VGND VGND VPWR VPWR _07858_/C sky130_fd_sc_hd__xnor2_4
XFILLER_44_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07769_ _07764_/A _07764_/B _07764_/C VGND VGND VPWR VPWR _07778_/B sky130_fd_sc_hd__a21o_1
XFILLER_112_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_36_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _13265_/CLK sky130_fd_sc_hd__clkbuf_16
X_09508_ _13605_/Q _13606_/Q _13607_/Q _13608_/Q _09562_/B VGND VGND VPWR VPWR _09508_/Y
+ sky130_fd_sc_hd__o41ai_4
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10780_ _10780_/A VGND VGND VPWR VPWR _13053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09439_ _09440_/B _09440_/C _13600_/Q VGND VGND VPWR VPWR _09448_/C sky130_fd_sc_hd__a21oi_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12450_ _14657_/Q _14514_/Q _12450_/S VGND VGND VPWR VPWR _12451_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11401_ _13724_/Q _11405_/B VGND VGND VPWR VPWR _11402_/A sky130_fd_sc_hd__and2_1
X_12381_ _12381_/A VGND VGND VPWR VPWR _14612_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_80 _12019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 _13094_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14120_ _14159_/CLK hold429/X VGND VGND VPWR VPWR _14120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11332_ _11332_/A VGND VGND VPWR VPWR _13770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14051_ _14703_/CLK _14051_/D VGND VGND VPWR VPWR _14051_/Q sky130_fd_sc_hd__dfxtp_1
X_11263_ _10944_/A _11260_/Y _11262_/Y _10929_/A VGND VGND VPWR VPWR _11264_/B sky130_fd_sc_hd__a211o_1
XFILLER_106_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13002_ _13525_/CLK _13002_/D hold1/X VGND VGND VPWR VPWR _13002_/Q sky130_fd_sc_hd__dfrtp_1
X_10214_ _14096_/Q _14080_/Q _14384_/D VGND VGND VPWR VPWR _10215_/A sky130_fd_sc_hd__mux2_1
X_11194_ _11242_/A _11194_/B VGND VGND VPWR VPWR _11194_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10145_ _14283_/D _10144_/X _14294_/D VGND VGND VPWR VPWR _10146_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10076_ _10076_/A VGND VGND VPWR VPWR _13887_/D sky130_fd_sc_hd__clkbuf_1
X_13904_ _14693_/CLK _13904_/D VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__dfxtp_1
XFILLER_75_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13835_ _14720_/CLK _13835_/D VGND VGND VPWR VPWR _13835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _13294_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13766_ _14714_/CLK _13766_/D VGND VGND VPWR VPWR _13766_/Q sky130_fd_sc_hd__dfxtp_1
X_10978_ _11037_/A _10978_/B VGND VGND VPWR VPWR _10978_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12717_ _13596_/CLK _12717_/D VGND VGND VPWR VPWR hold455/A sky130_fd_sc_hd__dfxtp_1
X_13697_ _13811_/CLK _13697_/D repeater57/X VGND VGND VPWR VPWR _13697_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_30_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12648_ _14743_/Q _12567_/X _12647_/X _12609_/X VGND VGND VPWR VPWR _14748_/D sky130_fd_sc_hd__o211a_1
XFILLER_62_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12579_ _12609_/A VGND VGND VPWR VPWR _12641_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14318_ _14726_/CLK _14318_/D VGND VGND VPWR VPWR _14318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold306 hold306/A VGND VGND VPWR VPWR hold306/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold317 hold317/A VGND VGND VPWR VPWR hold317/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold328 hold328/A VGND VGND VPWR VPWR hold328/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold339 hold339/A VGND VGND VPWR VPWR hold339/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_14249_ _14251_/CLK _14249_/D VGND VGND VPWR VPWR _14249_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08810_ _09006_/S VGND VGND VPWR VPWR _11268_/A sky130_fd_sc_hd__clkbuf_2
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09790_ _13677_/Q _09790_/B _09836_/D VGND VGND VPWR VPWR _09792_/A sky130_fd_sc_hd__and3_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _08741_/A _08741_/B _08741_/C _08739_/C VGND VGND VPWR VPWR _08742_/B sky130_fd_sc_hd__or4b_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05953_ _06161_/A VGND VGND VPWR VPWR _06309_/S sky130_fd_sc_hd__inv_2
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08672_ _09524_/B VGND VGND VPWR VPWR _09518_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_81_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07623_ _13113_/Q VGND VGND VPWR VPWR _07723_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_18_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _14098_/CLK sky130_fd_sc_hd__clkbuf_16
X_07554_ _07495_/X _07556_/B _07553_/Y _07499_/X VGND VGND VPWR VPWR _13157_/D sky130_fd_sc_hd__a31o_1
XFILLER_34_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06505_ _12885_/Q _06505_/B VGND VGND VPWR VPWR _06516_/A sky130_fd_sc_hd__nor2_1
XFILLER_50_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07485_ _07488_/A _07504_/B VGND VGND VPWR VPWR _07485_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09224_ _09242_/A _09223_/B _07524_/X VGND VGND VPWR VPWR _09224_/X sky130_fd_sc_hd__a21o_1
X_06436_ _06436_/A _06436_/B VGND VGND VPWR VPWR _06437_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06367_ _06365_/Y _06366_/X _14429_/D VGND VGND VPWR VPWR _06368_/A sky130_fd_sc_hd__mux2_1
X_09155_ _09156_/A _09156_/B _09156_/C VGND VGND VPWR VPWR _09155_/X sky130_fd_sc_hd__a21o_1
XFILLER_148_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08106_ _14012_/Q _14010_/Q _14008_/Q _14006_/Q _13424_/Q _08143_/A VGND VGND VPWR
+ VPWR _08209_/B sky130_fd_sc_hd__mux4_2
XFILLER_163_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06298_ _06298_/A VGND VGND VPWR VPWR _14209_/D sky130_fd_sc_hd__clkbuf_1
X_09086_ _13524_/Q _09086_/B _09086_/C VGND VGND VPWR VPWR _09089_/A sky130_fd_sc_hd__and3_1
XFILLER_163_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08037_ _08037_/A VGND VGND VPWR VPWR _12677_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09988_ _09987_/X _09984_/X _10596_/B VGND VGND VPWR VPWR _09989_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08939_ _08939_/A _08939_/B VGND VGND VPWR VPWR _08940_/B sky130_fd_sc_hd__nand2_1
XFILLER_123_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11950_ _14694_/Q VGND VGND VPWR VPWR _11950_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10901_ _10901_/A _10900_/Y VGND VGND VPWR VPWR _10901_/X sky130_fd_sc_hd__or2b_1
XFILLER_72_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11881_ _11881_/A VGND VGND VPWR VPWR _14237_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13620_ _13622_/CLK _13620_/D repeater57/X VGND VGND VPWR VPWR _13620_/Q sky130_fd_sc_hd__dfrtp_1
X_10832_ _10876_/A VGND VGND VPWR VPWR _10841_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13551_ _13552_/CLK _13551_/D _12609_/A VGND VGND VPWR VPWR _13551_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10763_ _10763_/A VGND VGND VPWR VPWR _13045_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12502_ _12502_/A _12502_/B input19/X VGND VGND VPWR VPWR _12503_/A sky130_fd_sc_hd__and3_1
Xrepeater59 hold1/X VGND VGND VPWR VPWR repeater59/X sky130_fd_sc_hd__buf_12
X_13482_ _13702_/CLK hold265/X VGND VGND VPWR VPWR _13482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10694_ _12883_/Q _10698_/B VGND VGND VPWR VPWR _10695_/A sky130_fd_sc_hd__and2_1
XFILLER_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12433_ _14649_/Q _14695_/Q _12439_/S VGND VGND VPWR VPWR _12434_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12364_ _14605_/Q _11981_/X _12364_/S VGND VGND VPWR VPWR _12365_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14103_ _14410_/CLK _14103_/D VGND VGND VPWR VPWR _14103_/Q sky130_fd_sc_hd__dfxtp_1
X_11315_ _13765_/Q _11313_/X _11327_/S VGND VGND VPWR VPWR _11316_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12295_ _12295_/A VGND VGND VPWR VPWR _14563_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14034_ _14724_/CLK _14034_/D VGND VGND VPWR VPWR _14034_/Q sky130_fd_sc_hd__dfxtp_1
X_11246_ _11246_/A _10960_/A VGND VGND VPWR VPWR _11246_/X sky130_fd_sc_hd__or2b_1
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11177_ _11177_/A _11177_/B VGND VGND VPWR VPWR _11177_/Y sky130_fd_sc_hd__nor2_1
X_10128_ _10128_/A VGND VGND VPWR VPWR _14178_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10059_ _10059_/A VGND VGND VPWR VPWR _14043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13818_ _14636_/CLK _13818_/D VGND VGND VPWR VPWR hold220/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13749_ _14588_/CLK _14583_/Q VGND VGND VPWR VPWR _13749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07270_ _07428_/A _07267_/X _07269_/X VGND VGND VPWR VPWR _07270_/X sky130_fd_sc_hd__a21o_1
X_06221_ _14395_/Q _14387_/Q _10197_/A VGND VGND VPWR VPWR _10626_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06152_ _14182_/Q _14174_/Q _06289_/S VGND VGND VPWR VPWR _06152_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold103 hold103/A VGND VGND VPWR VPWR hold103/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold114 hold114/A VGND VGND VPWR VPWR hold114/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_105_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06083_ _10606_/A _06082_/X _10034_/S VGND VGND VPWR VPWR _06084_/A sky130_fd_sc_hd__mux2_1
Xhold125 hold125/A VGND VGND VPWR VPWR hold125/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold136 hold136/A VGND VGND VPWR VPWR hold136/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_145_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _13314_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_160_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold147 hold147/A VGND VGND VPWR VPWR hold147/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold158 hold158/A VGND VGND VPWR VPWR hold158/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09911_ _13481_/Q _13670_/Q _09913_/S VGND VGND VPWR VPWR _09912_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold169 hold169/A VGND VGND VPWR VPWR hold169/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_125_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09842_ _09842_/A _09842_/B VGND VGND VPWR VPWR _09842_/Y sky130_fd_sc_hd__xnor2_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09773_ _09781_/A _09773_/B VGND VGND VPWR VPWR _09773_/Y sky130_fd_sc_hd__xnor2_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06985_ _13026_/Q _08002_/B VGND VGND VPWR VPWR _06986_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _08724_/A _08724_/B VGND VGND VPWR VPWR _08741_/B sky130_fd_sc_hd__nand2_1
X_05936_ _05923_/X _05924_/X _05928_/X _05935_/Y VGND VGND VPWR VPWR _05937_/B sky130_fd_sc_hd__a31o_1
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08655_ _08665_/A _09464_/B VGND VGND VPWR VPWR _08655_/X sky130_fd_sc_hd__and2_1
XFILLER_15_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ _07606_/A VGND VGND VPWR VPWR _13655_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08586_ _08591_/A _09424_/C _13444_/Q VGND VGND VPWR VPWR _08621_/A sky130_fd_sc_hd__a21oi_1
X_07537_ _07548_/A _07547_/A VGND VGND VPWR VPWR _07537_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07468_ _09237_/B VGND VGND VPWR VPWR _09258_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09207_ _13541_/Q _09207_/B VGND VGND VPWR VPWR _09208_/B sky130_fd_sc_hd__or2_1
X_06419_ _12878_/Q _06423_/B VGND VGND VPWR VPWR _06436_/A sky130_fd_sc_hd__or2_2
XFILLER_10_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07399_ _09125_/A VGND VGND VPWR VPWR _07399_/X sky130_fd_sc_hd__buf_2
XFILLER_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09138_ _09136_/X _09137_/Y _07365_/X _07326_/X VGND VGND VPWR VPWR _13531_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_136_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09069_ _13232_/Q _13461_/Q _09075_/S VGND VGND VPWR VPWR _09070_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11100_ _14024_/Q _13990_/Q _13830_/Q _14542_/Q _11081_/X _11082_/X VGND VGND VPWR
+ VPWR _11101_/A sky130_fd_sc_hd__mux4_1
XFILLER_78_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12080_ _12080_/A VGND VGND VPWR VPWR _14457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11031_ _10991_/X _11028_/X _11030_/X _11015_/X VGND VGND VPWR VPWR _11031_/X sky130_fd_sc_hd__o211a_1
XFILLER_1_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12982_ _13274_/CLK hold260/X VGND VGND VPWR VPWR _12982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14721_ _14721_/CLK _14721_/D VGND VGND VPWR VPWR _14721_/Q sky130_fd_sc_hd__dfxtp_1
X_11933_ _11933_/A VGND VGND VPWR VPWR _14272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14652_ _14652_/CLK _14652_/D VGND VGND VPWR VPWR _14652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ _14230_/Q _11478_/X _11864_/S VGND VGND VPWR VPWR _11865_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _13604_/CLK _13603_/D repeater56/X VGND VGND VPWR VPWR _13603_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _10815_/A VGND VGND VPWR VPWR _13069_/D sky130_fd_sc_hd__clkbuf_1
X_14583_ _14702_/CLK _14583_/D VGND VGND VPWR VPWR _14583_/Q sky130_fd_sc_hd__dfxtp_1
X_11795_ _13569_/Q _11795_/B VGND VGND VPWR VPWR _11796_/A sky130_fd_sc_hd__and2_1
XFILLER_41_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13534_ _13534_/CLK _13534_/D _12609_/A VGND VGND VPWR VPWR _13534_/Q sky130_fd_sc_hd__dfrtp_1
X_10746_ _12907_/Q _10748_/B VGND VGND VPWR VPWR _10747_/A sky130_fd_sc_hd__and2_1
X_13465_ _13622_/CLK _13465_/D repeater57/X VGND VGND VPWR VPWR _13465_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_159_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10677_ _13031_/D VGND VGND VPWR VPWR _10748_/B sky130_fd_sc_hd__buf_2
X_12416_ _12418_/A _12418_/B input3/X VGND VGND VPWR VPWR _12417_/A sky130_fd_sc_hd__and3_1
X_13396_ _13596_/CLK hold475/X VGND VGND VPWR VPWR _13396_/Q sky130_fd_sc_hd__dfxtp_1
X_12347_ _14597_/Q _11956_/X _12353_/S VGND VGND VPWR VPWR _12348_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12278_ _11375_/X _14554_/Q _12278_/S VGND VGND VPWR VPWR _12279_/A sky130_fd_sc_hd__mux2_1
X_14017_ _14707_/CLK _14017_/D VGND VGND VPWR VPWR _14017_/Q sky130_fd_sc_hd__dfxtp_1
X_11229_ _11240_/A _11229_/B VGND VGND VPWR VPWR _11229_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06770_ _06770_/A _06786_/B _06770_/C VGND VGND VPWR VPWR _07853_/B sky130_fd_sc_hd__nand3_1
XFILLER_36_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08440_ _09370_/B _08440_/B VGND VGND VPWR VPWR _13435_/D sky130_fd_sc_hd__xnor2_1
XFILLER_90_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08371_ _13083_/Q _13364_/Q _08373_/S VGND VGND VPWR VPWR _08372_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07322_ _07322_/A _07322_/B VGND VGND VPWR VPWR _07322_/X sky130_fd_sc_hd__xor2_1
XFILLER_31_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07253_ _13132_/Q _07261_/B _09086_/C VGND VGND VPWR VPWR _07255_/A sky130_fd_sc_hd__and3_1
XFILLER_164_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06204_ _06203_/X _06200_/X _10193_/A VGND VGND VPWR VPWR _06205_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07184_ _07209_/A _07184_/B VGND VGND VPWR VPWR _07184_/X sky130_fd_sc_hd__xor2_1
X_06135_ _06135_/A VGND VGND VPWR VPWR _14152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06066_ _13974_/Q _13972_/Q _10020_/A VGND VGND VPWR VPWR _06066_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09825_ _09821_/B _09824_/X _09834_/S VGND VGND VPWR VPWR _09826_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09756_ _09673_/X _09700_/X _09704_/B _09718_/Y VGND VGND VPWR VPWR _09758_/B sky130_fd_sc_hd__o22a_1
X_06968_ _06968_/A _06968_/B VGND VGND VPWR VPWR _06973_/C sky130_fd_sc_hd__nand2_1
XFILLER_86_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08707_ _13454_/Q _08730_/B VGND VGND VPWR VPWR _08714_/D sky130_fd_sc_hd__xnor2_1
X_05919_ _13726_/Q _13727_/Q _13728_/Q _13733_/Q VGND VGND VPWR VPWR _05920_/D sky130_fd_sc_hd__or4_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _09731_/A _14211_/Q VGND VGND VPWR VPWR _09687_/X sky130_fd_sc_hd__and2b_1
X_06899_ _06899_/A VGND VGND VPWR VPWR _06899_/Y sky130_fd_sc_hd__inv_2
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _09457_/B _09457_/C _13448_/Q VGND VGND VPWR VPWR _08653_/A sky130_fd_sc_hd__a21oi_1
XFILLER_27_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _09414_/B _09414_/C VGND VGND VPWR VPWR _08570_/A sky130_fd_sc_hd__and2_1
X_10600_ _10600_/A VGND VGND VPWR VPWR _13753_/D sky130_fd_sc_hd__inv_2
X_11580_ _11580_/A VGND VGND VPWR VPWR _13871_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10531_ _12991_/D _10531_/B VGND VGND VPWR VPWR _10534_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13250_ _13366_/CLK hold519/X VGND VGND VPWR VPWR hold504/A sky130_fd_sc_hd__dfxtp_1
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10462_ _10462_/A _10462_/B VGND VGND VPWR VPWR _10463_/B sky130_fd_sc_hd__xnor2_1
XFILLER_129_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12201_ _12201_/A VGND VGND VPWR VPWR _14511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13181_ _13434_/CLK _13181_/D VGND VGND VPWR VPWR hold353/A sky130_fd_sc_hd__dfxtp_1
X_10393_ _10393_/A _10393_/B VGND VGND VPWR VPWR _10394_/B sky130_fd_sc_hd__nor2_1
XFILLER_136_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12132_ _12132_/A VGND VGND VPWR VPWR _14480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12063_ _11310_/X _14450_/Q _12063_/S VGND VGND VPWR VPWR _12064_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11014_ _11014_/A _11013_/X VGND VGND VPWR VPWR _11014_/X sky130_fd_sc_hd__or2b_1
XFILLER_77_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12965_ _13265_/CLK hold391/X VGND VGND VPWR VPWR _12965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14704_ _14704_/CLK _14704_/D VGND VGND VPWR VPWR _14704_/Q sky130_fd_sc_hd__dfxtp_1
X_11916_ _14265_/Q _11475_/X _11918_/S VGND VGND VPWR VPWR _11917_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12896_ _12970_/CLK _12896_/D repeater59/X VGND VGND VPWR VPWR _12896_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _14636_/CLK _14635_/D VGND VGND VPWR VPWR hold322/A sky130_fd_sc_hd__dfxtp_1
X_11847_ _14222_/Q _11453_/X _11853_/S VGND VGND VPWR VPWR _11848_/A sky130_fd_sc_hd__mux2_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _14605_/CLK _14566_/D VGND VGND VPWR VPWR _14566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11778_ _13561_/Q _11784_/B VGND VGND VPWR VPWR _11779_/A sky130_fd_sc_hd__and2_1
XFILLER_158_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13517_ _13520_/CLK _13517_/D VGND VGND VPWR VPWR _13517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10729_ _12899_/Q _10731_/B VGND VGND VPWR VPWR _10730_/A sky130_fd_sc_hd__and2_1
X_14497_ _14605_/CLK _14497_/D VGND VGND VPWR VPWR _14497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13448_ _13602_/CLK _13448_/D repeater56/X VGND VGND VPWR VPWR _13448_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_155_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13379_ _14333_/CLK _13379_/D _12609_/A VGND VGND VPWR VPWR _13379_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07940_ _07940_/A VGND VGND VPWR VPWR _07940_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07871_ _07885_/A _07885_/C VGND VGND VPWR VPWR _07884_/C sky130_fd_sc_hd__nor2_1
X_09610_ _09610_/A VGND VGND VPWR VPWR _12819_/D sky130_fd_sc_hd__clkbuf_1
X_06822_ _06665_/X _06819_/X _06820_/Y _06821_/X VGND VGND VPWR VPWR _13009_/D sky130_fd_sc_hd__a31o_1
XFILLER_83_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09541_ _09539_/Y _09540_/X _09493_/X VGND VGND VPWR VPWR _13613_/D sky130_fd_sc_hd__a21o_1
X_06753_ _06753_/A _06753_/B _06753_/C VGND VGND VPWR VPWR _06786_/B sky130_fd_sc_hd__and3_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09472_ _13604_/Q _09472_/B VGND VGND VPWR VPWR _09473_/B sky130_fd_sc_hd__nor2_1
X_06684_ _06895_/A VGND VGND VPWR VPWR _06859_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08423_ _13249_/Q _13433_/Q VGND VGND VPWR VPWR _09002_/A sky130_fd_sc_hd__xor2_2
XFILLER_24_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08354_ _13075_/Q _13356_/Q _08362_/S VGND VGND VPWR VPWR _08355_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07305_ _07305_/A _07305_/B _07305_/C VGND VGND VPWR VPWR _07321_/B sky130_fd_sc_hd__or3_1
X_08285_ _08285_/A _08285_/B VGND VGND VPWR VPWR _08285_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_138_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07236_ _13131_/Q _08124_/A VGND VGND VPWR VPWR _07237_/B sky130_fd_sc_hd__nand2_1
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07167_ _07142_/A _07144_/B _07142_/B VGND VGND VPWR VPWR _07168_/A sky130_fd_sc_hd__o21ba_1
XFILLER_145_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06118_ _14207_/Q _14205_/Q _14209_/Q VGND VGND VPWR VPWR _06119_/B sky130_fd_sc_hd__mux2_1
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07098_ _07098_/A _07098_/B VGND VGND VPWR VPWR _07131_/A sky130_fd_sc_hd__xnor2_1
X_06049_ _13929_/Q _06049_/B VGND VGND VPWR VPWR _06057_/A sky130_fd_sc_hd__xnor2_2
XFILLER_87_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09808_ _09808_/A VGND VGND VPWR VPWR _13678_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09739_ _13672_/Q _09739_/B VGND VGND VPWR VPWR _09741_/A sky130_fd_sc_hd__xnor2_1
XFILLER_28_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12750_ _13702_/CLK _12750_/D VGND VGND VPWR VPWR hold168/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11701_/A VGND VGND VPWR VPWR _14032_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _13296_/CLK _12681_/D VGND VGND VPWR VPWR hold382/A sky130_fd_sc_hd__dfxtp_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14732_/CLK _14420_/D VGND VGND VPWR VPWR _14420_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _13992_/Q _11491_/X _11634_/S VGND VGND VPWR VPWR _11633_/A sky130_fd_sc_hd__mux2_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14351_ _14557_/CLK _14351_/D VGND VGND VPWR VPWR hold106/A sky130_fd_sc_hd__dfxtp_1
X_11563_ _13640_/Q _11563_/B VGND VGND VPWR VPWR _11564_/A sky130_fd_sc_hd__and2_1
XFILLER_156_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13302_ _13574_/CLK hold24/X VGND VGND VPWR VPWR _13302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10514_ _10514_/A VGND VGND VPWR VPWR _14433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14282_ _14294_/CLK _14282_/D VGND VGND VPWR VPWR _14282_/Q sky130_fd_sc_hd__dfxtp_1
X_11494_ _14519_/Q VGND VGND VPWR VPWR _11494_/X sky130_fd_sc_hd__buf_2
X_13233_ _13617_/CLK hold449/X VGND VGND VPWR VPWR _13233_/Q sky130_fd_sc_hd__dfxtp_1
X_10445_ hold64/A VGND VGND VPWR VPWR _10495_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13164_ _13562_/CLK hold23/X VGND VGND VPWR VPWR _13468_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_152_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10376_ _10376_/A _10423_/A _10376_/C VGND VGND VPWR VPWR _10396_/A sky130_fd_sc_hd__and3_1
X_12115_ _14473_/Q _11978_/X _12117_/S VGND VGND VPWR VPWR _12116_/A sky130_fd_sc_hd__mux2_1
X_13095_ _13587_/CLK hold298/X VGND VGND VPWR VPWR _13095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12046_ _11285_/X _14442_/Q _12052_/S VGND VGND VPWR VPWR _12047_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13997_ _14721_/CLK _13997_/D VGND VGND VPWR VPWR _13997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12948_ _13314_/CLK _12948_/D VGND VGND VPWR VPWR hold214/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ _12881_/CLK _12879_/D hold1/X VGND VGND VPWR VPWR _12879_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14618_ _14619_/CLK _14618_/D VGND VGND VPWR VPWR _14618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14549_ _14721_/CLK _14549_/D VGND VGND VPWR VPWR _14549_/Q sky130_fd_sc_hd__dfxtp_1
X_08070_ _08070_/A VGND VGND VPWR VPWR _12695_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07021_ _10339_/A hold131/A VGND VGND VPWR VPWR _07218_/S sky130_fd_sc_hd__xor2_4
XFILLER_115_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08972_ _08997_/A _08972_/B VGND VGND VPWR VPWR _08972_/X sky130_fd_sc_hd__xor2_1
XFILLER_142_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07923_ _07923_/A _07923_/B VGND VGND VPWR VPWR _07949_/A sky130_fd_sc_hd__nand2_1
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_57_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07854_ _07853_/B _07853_/C _13260_/Q VGND VGND VPWR VPWR _07885_/B sky130_fd_sc_hd__a21oi_1
XFILLER_56_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06805_ _06825_/A _06806_/B VGND VGND VPWR VPWR _06820_/B sky130_fd_sc_hd__or2_1
X_07785_ _07745_/C _07785_/B _07785_/C VGND VGND VPWR VPWR _07789_/A sky130_fd_sc_hd__and3b_1
XFILLER_72_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09524_ _13611_/Q _09524_/B VGND VGND VPWR VPWR _09532_/A sky130_fd_sc_hd__and2_1
X_06736_ _06736_/A _06736_/B VGND VGND VPWR VPWR _06753_/B sky130_fd_sc_hd__and2_2
XFILLER_64_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09455_ _09455_/A _09455_/B _09455_/C VGND VGND VPWR VPWR _09455_/Y sky130_fd_sc_hd__nand3_1
X_06667_ _13036_/Q _13352_/Q _06705_/S VGND VGND VPWR VPWR _06852_/B sky130_fd_sc_hd__mux2_1
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08406_ _13099_/Q _13380_/Q _08406_/S VGND VGND VPWR VPWR _08407_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09386_ _09388_/B _09385_/Y _09404_/S VGND VGND VPWR VPWR _09387_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06598_ _12898_/Q _12899_/Q _06598_/C _06598_/D VGND VGND VPWR VPWR _06607_/D sky130_fd_sc_hd__and4_1
XFILLER_101_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08337_ _08331_/A _13382_/Q _08331_/B _13383_/Q VGND VGND VPWR VPWR _08338_/B sky130_fd_sc_hd__a31o_1
XFILLER_131_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08268_ _09125_/A _08268_/B VGND VGND VPWR VPWR _08268_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07219_ _07219_/A VGND VGND VPWR VPWR _13353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08199_ _08199_/A _08199_/B _08199_/C VGND VGND VPWR VPWR _08201_/B sky130_fd_sc_hd__and3_1
XFILLER_134_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10230_ _10230_/A VGND VGND VPWR VPWR _10230_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10161_ _14288_/D _10160_/X _14293_/D VGND VGND VPWR VPWR _10161_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10092_ _10085_/X _13908_/D _10092_/S VGND VGND VPWR VPWR _10092_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13920_ _14042_/CLK _13920_/D VGND VGND VPWR VPWR _13920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13851_ _14180_/CLK _13851_/D VGND VGND VPWR VPWR _13851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12802_ _14275_/CLK _12802_/D VGND VGND VPWR VPWR hold164/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13782_ _14647_/CLK _13814_/Q VGND VGND VPWR VPWR _13782_/Q sky130_fd_sc_hd__dfxtp_1
X_10994_ _11163_/A VGND VGND VPWR VPWR _10995_/A sky130_fd_sc_hd__buf_2
XFILLER_55_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12733_ _14696_/CLK _12733_/D VGND VGND VPWR VPWR hold379/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12664_ _14702_/CLK _12664_/D VGND VGND VPWR VPWR _13245_/D sky130_fd_sc_hd__dfxtp_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _14410_/CLK _14403_/D VGND VGND VPWR VPWR _14403_/Q sky130_fd_sc_hd__dfxtp_1
X_11615_ _13984_/Q _11465_/X _11623_/S VGND VGND VPWR VPWR _11616_/A sky130_fd_sc_hd__mux2_1
X_12595_ _12595_/A VGND VGND VPWR VPWR _14728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14334_ _14697_/CLK hold29/X VGND VGND VPWR VPWR _14334_/Q sky130_fd_sc_hd__dfxtp_1
X_11546_ _13632_/Q _11552_/B VGND VGND VPWR VPWR _11547_/A sky130_fd_sc_hd__and2_1
XFILLER_128_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14265_ _14656_/CLK _14265_/D VGND VGND VPWR VPWR _14265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11477_ _11477_/A VGND VGND VPWR VPWR _13827_/D sky130_fd_sc_hd__clkbuf_1
X_13216_ _13423_/CLK hold367/X VGND VGND VPWR VPWR _13216_/Q sky130_fd_sc_hd__dfxtp_1
X_10428_ _10428_/A VGND VGND VPWR VPWR _14219_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14196_ _14196_/CLK _14196_/D VGND VGND VPWR VPWR _14196_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _13555_/CLK _13147_/D _12609_/A VGND VGND VPWR VPWR _13147_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _13782_/Q _10359_/B VGND VGND VPWR VPWR _12988_/D sky130_fd_sc_hd__xnor2_1
XFILLER_152_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _13528_/CLK hold305/X VGND VGND VPWR VPWR _13078_/Q sky130_fd_sc_hd__dfxtp_1
X_12029_ _12029_/A VGND VGND VPWR VPWR _14323_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07570_ _08124_/A VGND VGND VPWR VPWR _07570_/X sky130_fd_sc_hd__buf_2
XFILLER_65_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06521_ _06514_/B _06520_/Y _06530_/S VGND VGND VPWR VPWR _06522_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09240_ _09125_/X _09239_/Y _07486_/X VGND VGND VPWR VPWR _13546_/D sky130_fd_sc_hd__a21o_1
X_06452_ _06452_/A _06452_/B VGND VGND VPWR VPWR _06452_/X sky130_fd_sc_hd__xor2_1
XFILLER_33_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09171_ _09177_/A _09177_/B VGND VGND VPWR VPWR _09172_/B sky130_fd_sc_hd__and2_1
X_06383_ _13107_/D VGND VGND VPWR VPWR _06455_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08122_ _08122_/A _08121_/X VGND VGND VPWR VPWR _08123_/B sky130_fd_sc_hd__or2b_1
XFILLER_147_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14755__66 VGND VGND VPWR VPWR _14755__66/HI data_o[29] sky130_fd_sc_hd__conb_1
XFILLER_135_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08053_ _10803_/A VGND VGND VPWR VPWR _08062_/S sky130_fd_sc_hd__buf_2
XFILLER_116_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07004_ _13029_/Q _08020_/B VGND VGND VPWR VPWR _07004_/X sky130_fd_sc_hd__or2_1
XFILLER_116_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08955_ _08930_/A _08932_/B _08930_/B VGND VGND VPWR VPWR _08956_/A sky130_fd_sc_hd__o21ba_1
XFILLER_69_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07906_ _07916_/A _07906_/B VGND VGND VPWR VPWR _07914_/B sky130_fd_sc_hd__or2_1
X_08886_ _08886_/A _08886_/B VGND VGND VPWR VPWR _08919_/A sky130_fd_sc_hd__xnor2_1
XFILLER_57_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07837_ _07811_/X _07835_/Y _07836_/X _06733_/X VGND VGND VPWR VPWR _13257_/D sky130_fd_sc_hd__a31o_1
XFILLER_72_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07768_ _07768_/A VGND VGND VPWR VPWR _13662_/D sky130_fd_sc_hd__clkbuf_1
X_09507_ _09502_/X _09504_/X _09505_/Y _09506_/X VGND VGND VPWR VPWR _13608_/D sky130_fd_sc_hd__a31o_1
X_06719_ _06719_/A VGND VGND VPWR VPWR _06770_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_07699_ _13115_/Q VGND VGND VPWR VPWR _07772_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09438_ _13599_/Q _09438_/B VGND VGND VPWR VPWR _09443_/A sky130_fd_sc_hd__nand2_1
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09369_ _09369_/A _09368_/X VGND VGND VPWR VPWR _09371_/A sky130_fd_sc_hd__or2b_1
XFILLER_138_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11400_ _11400_/A VGND VGND VPWR VPWR _13792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12380_ _14612_/Q _12004_/X _12386_/S VGND VGND VPWR VPWR _12381_/A sky130_fd_sc_hd__mux2_1
XANTENNA_70 _13551_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_81 _12022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11331_ _13770_/Q _11329_/X _11355_/S VGND VGND VPWR VPWR _11332_/A sky130_fd_sc_hd__mux2_1
XANTENNA_92 _13031_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14050_ _14050_/CLK _14050_/D VGND VGND VPWR VPWR _14050_/Q sky130_fd_sc_hd__dfxtp_1
X_11262_ _11262_/A _11262_/B VGND VGND VPWR VPWR _11262_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13001_ _13525_/CLK _13001_/D hold1/X VGND VGND VPWR VPWR _13001_/Q sky130_fd_sc_hd__dfrtp_1
X_10213_ _10213_/A VGND VGND VPWR VPWR _14394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11193_ _11159_/X _11189_/Y _11192_/Y _11166_/X VGND VGND VPWR VPWR _11194_/B sky130_fd_sc_hd__a211o_1
XFILLER_106_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10144_ _14152_/Q _10143_/X _10147_/A VGND VGND VPWR VPWR _10144_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_2_0_0_clk clkbuf_2_1_0_clk/A VGND VGND VPWR VPWR clkbuf_3_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10075_ _14046_/D _10074_/X _14048_/D VGND VGND VPWR VPWR _10076_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13903_ _14210_/CLK _13903_/D VGND VGND VPWR VPWR hold148/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13834_ _14275_/CLK _13834_/D VGND VGND VPWR VPWR _13834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13765_ _14713_/CLK _13765_/D VGND VGND VPWR VPWR _13765_/Q sky130_fd_sc_hd__dfxtp_1
X_10977_ _10932_/X _10972_/Y _10976_/Y _10946_/X VGND VGND VPWR VPWR _10978_/B sky130_fd_sc_hd__a211o_1
XFILLER_31_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12716_ _13596_/CLK _12716_/D VGND VGND VPWR VPWR hold415/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13696_ _13811_/CLK _13696_/D repeater57/X VGND VGND VPWR VPWR _13696_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12647_ _12647_/A _12649_/B VGND VGND VPWR VPWR _12647_/X sky130_fd_sc_hd__or2_1
XFILLER_12_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12578_ _12567_/X _12572_/Y _12577_/X _10901_/X VGND VGND VPWR VPWR _12578_/X sky130_fd_sc_hd__o31a_1
XFILLER_144_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14317_ _14619_/CLK _14317_/D VGND VGND VPWR VPWR _14317_/Q sky130_fd_sc_hd__dfxtp_1
X_11529_ _13625_/Q _11529_/B VGND VGND VPWR VPWR _11530_/A sky130_fd_sc_hd__and2_1
XFILLER_156_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold307 hold307/A VGND VGND VPWR VPWR hold307/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold318 hold318/A VGND VGND VPWR VPWR hold318/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold329 hold329/A VGND VGND VPWR VPWR hold329/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_14248_ _14250_/CLK _14248_/D VGND VGND VPWR VPWR _14248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14179_ _14179_/CLK _14179_/D VGND VGND VPWR VPWR _14179_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _08706_/X _08738_/Y _08739_/X _08696_/X VGND VGND VPWR VPWR _13458_/D sky130_fd_sc_hd__a31o_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05952_ _05952_/A _05952_/B VGND VGND VPWR VPWR _06161_/A sky130_fd_sc_hd__nor2_1
XFILLER_38_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08671_ _08671_/A _08671_/B _08671_/C VGND VGND VPWR VPWR _09524_/B sky130_fd_sc_hd__and3_2
XFILLER_54_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07622_ _07622_/A _07747_/A VGND VGND VPWR VPWR _07641_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07553_ _07559_/A _07553_/B _07553_/C VGND VGND VPWR VPWR _07553_/Y sky130_fd_sc_hd__nand3_1
XFILLER_81_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06504_ _12885_/Q _06504_/B _06554_/C VGND VGND VPWR VPWR _06506_/A sky130_fd_sc_hd__and3_1
XFILLER_22_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07484_ _07488_/A _07504_/B VGND VGND VPWR VPWR _07484_/X sky130_fd_sc_hd__or2_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09223_ _09242_/A _09223_/B VGND VGND VPWR VPWR _09226_/B sky130_fd_sc_hd__nor2_1
X_06435_ _12876_/Q _06391_/A _06399_/B _06434_/X _06397_/X VGND VGND VPWR VPWR _06436_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09154_ _09159_/B _09159_/C VGND VGND VPWR VPWR _09156_/C sky130_fd_sc_hd__or2_1
X_06366_ _14645_/Q _14428_/D VGND VGND VPWR VPWR _06366_/X sky130_fd_sc_hd__and2_1
XFILLER_148_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08105_ _13425_/Q VGND VGND VPWR VPWR _08143_/A sky130_fd_sc_hd__clkbuf_2
X_09085_ _09088_/B _09085_/B VGND VGND VPWR VPWR _13523_/D sky130_fd_sc_hd__xnor2_1
X_06297_ _06295_/Y _06296_/X _14207_/D VGND VGND VPWR VPWR _06298_/A sky130_fd_sc_hd__mux2_1
X_08036_ _12956_/Q _13256_/Q _08040_/S VGND VGND VPWR VPWR _08037_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09987_ _14594_/Q _14592_/Q _13754_/Q VGND VGND VPWR VPWR _09987_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08938_ _08938_/A _08938_/B VGND VGND VPWR VPWR _08940_/A sky130_fd_sc_hd__xnor2_1
X_08869_ _08869_/A VGND VGND VPWR VPWR _14248_/D sky130_fd_sc_hd__clkbuf_1
X_10900_ _14749_/Q _14739_/Q VGND VGND VPWR VPWR _10900_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_17_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11880_ _14237_/Q _11501_/X _11886_/S VGND VGND VPWR VPWR _11881_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10831_ _10831_/A VGND VGND VPWR VPWR _10876_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13550_ _14530_/CLK _13550_/D _12609_/A VGND VGND VPWR VPWR _13550_/Q sky130_fd_sc_hd__dfrtp_4
X_10762_ _13003_/Q _10768_/B VGND VGND VPWR VPWR _10763_/A sky130_fd_sc_hd__and2_1
X_12501_ _12501_/A VGND VGND VPWR VPWR _14680_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13481_ _14250_/CLK hold183/X VGND VGND VPWR VPWR _13481_/Q sky130_fd_sc_hd__dfxtp_1
X_10693_ _10693_/A VGND VGND VPWR VPWR _12925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12432_ _12432_/A VGND VGND VPWR VPWR _14648_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12363_ _12363_/A VGND VGND VPWR VPWR _14604_/D sky130_fd_sc_hd__clkbuf_1
X_14102_ _14108_/CLK _14102_/D VGND VGND VPWR VPWR _14102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11314_ _11330_/A VGND VGND VPWR VPWR _11327_/S sky130_fd_sc_hd__buf_2
X_12294_ _14563_/Q _11968_/X _12302_/S VGND VGND VPWR VPWR _12295_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14033_ _14724_/CLK _14033_/D VGND VGND VPWR VPWR _14033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11245_ _14035_/Q _14001_/Q _13841_/Q _14553_/Q _10993_/A _10995_/A VGND VGND VPWR
+ VPWR _11246_/A sky130_fd_sc_hd__mux4_1
XFILLER_79_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11176_ _14273_/Q _14664_/Q _13771_/Q _14719_/Q _11162_/X _11163_/X VGND VGND VPWR
+ VPWR _11177_/B sky130_fd_sc_hd__mux4_1
XFILLER_121_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10127_ _13864_/Q _13848_/Q _14167_/D VGND VGND VPWR VPWR _10128_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10058_ _14039_/D _10057_/X _14050_/D VGND VGND VPWR VPWR _10059_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13817_ _14636_/CLK hold220/X VGND VGND VPWR VPWR hold211/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13748_ _14010_/CLK _13748_/D VGND VGND VPWR VPWR _13748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13679_ _13680_/CLK _13679_/D repeater56/X VGND VGND VPWR VPWR _13679_/Q sky130_fd_sc_hd__dfrtp_1
X_06220_ _06321_/S VGND VGND VPWR VPWR _10197_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_157_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06151_ _14178_/Q _14170_/Q _10110_/A VGND VGND VPWR VPWR _10616_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold104 hold104/A VGND VGND VPWR VPWR hold104/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_145_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold115 hold30/X VGND VGND VPWR VPWR hold115/X sky130_fd_sc_hd__clkbuf_1
X_06082_ _13950_/Q _13942_/Q _06256_/S VGND VGND VPWR VPWR _06082_/X sky130_fd_sc_hd__mux2_1
Xhold126 hold126/A VGND VGND VPWR VPWR hold126/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold137 hold137/A VGND VGND VPWR VPWR hold137/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold148 hold148/A VGND VGND VPWR VPWR hold148/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_160_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09910_ _09910_/A VGND VGND VPWR VPWR _12843_/D sky130_fd_sc_hd__clkbuf_1
Xhold159 hold159/A VGND VGND VPWR VPWR hold159/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09841_ _09840_/Y _09833_/B _09830_/A VGND VGND VPWR VPWR _09842_/B sky130_fd_sc_hd__a21oi_1
XFILLER_113_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09772_ _09753_/A _09753_/B _09763_/A _09771_/Y VGND VGND VPWR VPWR _09773_/B sky130_fd_sc_hd__o31ai_4
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06984_ _13026_/Q _08001_/B VGND VGND VPWR VPWR _06986_/A sky130_fd_sc_hd__and2_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _13456_/Q _09530_/B VGND VGND VPWR VPWR _08724_/B sky130_fd_sc_hd__or2_1
X_05935_ _05935_/A _05935_/B _05935_/C VGND VGND VPWR VPWR _05935_/Y sky130_fd_sc_hd__nor3_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08654_ _08654_/A _08654_/B VGND VGND VPWR VPWR _08664_/B sky130_fd_sc_hd__or2_1
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07605_ _11266_/B _07602_/Y _11266_/A VGND VGND VPWR VPWR _07606_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08585_ _13444_/Q _08591_/A _09424_/C VGND VGND VPWR VPWR _08587_/A sky130_fd_sc_hd__and3_1
XFILLER_156_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07536_ _13155_/Q _09257_/B VGND VGND VPWR VPWR _07547_/A sky130_fd_sc_hd__xor2_2
XFILLER_41_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07467_ _09212_/B VGND VGND VPWR VPWR _09237_/B sky130_fd_sc_hd__buf_2
XFILLER_22_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09206_ _13541_/Q _09206_/B VGND VGND VPWR VPWR _09214_/A sky130_fd_sc_hd__nand2_1
X_06418_ _06482_/A _06513_/B _06417_/X _06471_/A VGND VGND VPWR VPWR _06423_/B sky130_fd_sc_hd__o211a_1
X_07398_ _08303_/A VGND VGND VPWR VPWR _09125_/A sky130_fd_sc_hd__buf_2
XFILLER_5_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09137_ _09161_/A _09137_/B VGND VGND VPWR VPWR _09137_/Y sky130_fd_sc_hd__nor2_1
X_06349_ hold77/A _14401_/D _14402_/D _14405_/D VGND VGND VPWR VPWR _06350_/D sky130_fd_sc_hd__or4_1
XFILLER_135_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09068_ _09068_/A VGND VGND VPWR VPWR _12767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08019_ _06793_/A _08017_/X _08018_/Y _06930_/X VGND VGND VPWR VPWR _13282_/D sky130_fd_sc_hd__a31o_1
XFILLER_135_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11030_ _11030_/A _11013_/X VGND VGND VPWR VPWR _11030_/X sky130_fd_sc_hd__or2b_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12981_ _13314_/CLK hold214/X VGND VGND VPWR VPWR _12981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14720_ _14720_/CLK _14720_/D VGND VGND VPWR VPWR _14720_/Q sky130_fd_sc_hd__dfxtp_1
X_11932_ _14272_/Q _11497_/X _11940_/S VGND VGND VPWR VPWR _11933_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11863_ _11863_/A VGND VGND VPWR VPWR _14229_/D sky130_fd_sc_hd__clkbuf_1
X_14651_ _14652_/CLK _14651_/D VGND VGND VPWR VPWR _14651_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _13027_/Q _10818_/B VGND VGND VPWR VPWR _10815_/A sky130_fd_sc_hd__and2_1
X_13602_ _13602_/CLK _13602_/D repeater57/X VGND VGND VPWR VPWR _13602_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14582_ _14702_/CLK _14688_/Q VGND VGND VPWR VPWR hold101/A sky130_fd_sc_hd__dfxtp_1
X_11794_ _11794_/A VGND VGND VPWR VPWR _14090_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10745_ _10745_/A VGND VGND VPWR VPWR _12949_/D sky130_fd_sc_hd__clkbuf_1
X_13533_ _13534_/CLK _13533_/D _12609_/A VGND VGND VPWR VPWR _13533_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_158_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13464_ _13622_/CLK _13464_/D repeater57/X VGND VGND VPWR VPWR _13464_/Q sky130_fd_sc_hd__dfrtp_1
X_10676_ _14343_/Q _10671_/X _10675_/Y VGND VGND VPWR VPWR _12918_/D sky130_fd_sc_hd__o21a_1
XFILLER_71_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12415_ _12415_/A VGND VGND VPWR VPWR _14641_/D sky130_fd_sc_hd__clkbuf_1
X_13395_ _13596_/CLK hold377/X VGND VGND VPWR VPWR _13395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12346_ _12346_/A VGND VGND VPWR VPWR _14596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12277_ _12277_/A VGND VGND VPWR VPWR _14553_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14016_ _14707_/CLK _14016_/D VGND VGND VPWR VPWR _14016_/Q sky130_fd_sc_hd__dfxtp_1
X_11228_ _14277_/Q _14668_/Q _13775_/Q _14723_/Q _10914_/A _10918_/A VGND VGND VPWR
+ VPWR _11229_/B sky130_fd_sc_hd__mux4_1
X_11159_ _11190_/A VGND VGND VPWR VPWR _11159_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08370_ _08370_/A VGND VGND VPWR VPWR _12718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07321_ _07321_/A _07321_/B VGND VGND VPWR VPWR _07322_/B sky130_fd_sc_hd__and2_1
XFILLER_20_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07252_ _07461_/B _07249_/C _07249_/D _07461_/A VGND VGND VPWR VPWR _09086_/C sky130_fd_sc_hd__a22o_1
XFILLER_118_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06203_ _14422_/Q _14420_/Q _10194_/A VGND VGND VPWR VPWR _06203_/X sky130_fd_sc_hd__mux2_1
X_07183_ _07183_/A _07183_/B VGND VGND VPWR VPWR _07184_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06134_ _06133_/X _06130_/X _10106_/A VGND VGND VPWR VPWR _06135_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06065_ _06065_/A VGND VGND VPWR VPWR _13920_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09824_ _09824_/A _09824_/B VGND VGND VPWR VPWR _09824_/X sky130_fd_sc_hd__xor2_1
XFILLER_100_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06967_ _06967_/A _06967_/B VGND VGND VPWR VPWR _06968_/B sky130_fd_sc_hd__and2_1
XFILLER_101_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09755_ _09755_/A VGND VGND VPWR VPWR _13673_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08706_ _09502_/A VGND VGND VPWR VPWR _08706_/X sky130_fd_sc_hd__clkbuf_2
X_05918_ _13722_/Q _13723_/Q _13724_/Q _13725_/Q VGND VGND VPWR VPWR _05921_/C sky130_fd_sc_hd__or4_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09686_ _14220_/Q _09731_/A VGND VGND VPWR VPWR _09827_/B sky130_fd_sc_hd__and2_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06898_ _06874_/X _06888_/Y _06897_/X VGND VGND VPWR VPWR _13014_/D sky130_fd_sc_hd__a21o_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08637_ _13448_/Q _09457_/B _09457_/C VGND VGND VPWR VPWR _08644_/A sky130_fd_sc_hd__and3_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _08521_/A _08582_/B _08567_/C VGND VGND VPWR VPWR _09414_/C sky130_fd_sc_hd__a21o_1
X_07519_ _07519_/A _07515_/B VGND VGND VPWR VPWR _07519_/X sky130_fd_sc_hd__or2b_1
XFILLER_23_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08499_ _08481_/A _08477_/Y _08480_/B VGND VGND VPWR VPWR _08500_/B sky130_fd_sc_hd__o21a_1
X_10530_ _12991_/D _10537_/A VGND VGND VPWR VPWR _10547_/A sky130_fd_sc_hd__and2_1
XFILLER_127_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10461_ _10456_/X _10461_/B VGND VGND VPWR VPWR _10462_/B sky130_fd_sc_hd__and2b_1
XFILLER_136_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12200_ _14511_/Q _12022_/X _12202_/S VGND VGND VPWR VPWR _12201_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13180_ _13596_/CLK _13180_/D VGND VGND VPWR VPWR _13213_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_129_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10392_ _10393_/A _10393_/B VGND VGND VPWR VPWR _10407_/B sky130_fd_sc_hd__and2_1
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12131_ _14480_/Q _12000_/X _12139_/S VGND VGND VPWR VPWR _12132_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12062_ _12062_/A VGND VGND VPWR VPWR _14449_/D sky130_fd_sc_hd__clkbuf_1
Xhold490 hold13/X VGND VGND VPWR VPWR hold490/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_151_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11013_ _11155_/A VGND VGND VPWR VPWR _11013_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12964_ _13265_/CLK hold282/X VGND VGND VPWR VPWR _12964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14703_ _14703_/CLK _14703_/D VGND VGND VPWR VPWR _14703_/Q sky130_fd_sc_hd__dfxtp_1
X_11915_ _11915_/A VGND VGND VPWR VPWR _14264_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12895_ _12970_/CLK _12895_/D hold1/X VGND VGND VPWR VPWR _12895_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14634_ _14634_/CLK _14634_/D VGND VGND VPWR VPWR _14634_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _11846_/A VGND VGND VPWR VPWR _14221_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565_ _14605_/CLK _14565_/D VGND VGND VPWR VPWR _14565_/Q sky130_fd_sc_hd__dfxtp_1
X_11777_ _11777_/A VGND VGND VPWR VPWR _14082_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13516_ _13520_/CLK _13516_/D VGND VGND VPWR VPWR _13516_/Q sky130_fd_sc_hd__dfxtp_1
X_10728_ _10728_/A VGND VGND VPWR VPWR _12941_/D sky130_fd_sc_hd__clkbuf_1
X_14496_ _14712_/CLK _14496_/D VGND VGND VPWR VPWR _14496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10659_ _14337_/Q _14334_/Q _14338_/Q VGND VGND VPWR VPWR _10666_/C sky130_fd_sc_hd__and3_1
X_13447_ _13704_/CLK _13447_/D repeater56/X VGND VGND VPWR VPWR _13447_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13378_ _14696_/CLK _13378_/D _12609_/A VGND VGND VPWR VPWR _13378_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12329_ _12329_/A VGND VGND VPWR VPWR _14579_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07870_ _13262_/Q _07876_/B VGND VGND VPWR VPWR _07892_/B sky130_fd_sc_hd__xnor2_2
XFILLER_69_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06821_ _06871_/A _07878_/B _07878_/C VGND VGND VPWR VPWR _06821_/X sky130_fd_sc_hd__and3_1
XFILLER_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09540_ _09548_/A _09547_/A _08633_/A VGND VGND VPWR VPWR _09540_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06752_ _06745_/X _06863_/B _06751_/X _06736_/A VGND VGND VPWR VPWR _06753_/C sky130_fd_sc_hd__o211a_1
XFILLER_37_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09471_ _13604_/Q _09471_/B VGND VGND VPWR VPWR _09473_/A sky130_fd_sc_hd__and2_1
X_06683_ _13032_/Q VGND VGND VPWR VPWR _06895_/A sky130_fd_sc_hd__clkinv_2
XFILLER_24_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08422_ _08422_/A VGND VGND VPWR VPWR _12741_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08353_ _08397_/A VGND VGND VPWR VPWR _08362_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_11_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07304_ _07276_/A _07276_/B _07292_/Y _07290_/X VGND VGND VPWR VPWR _07305_/C sky130_fd_sc_hd__o211a_1
X_08284_ _08283_/Y _08276_/B _08273_/A VGND VGND VPWR VPWR _08285_/B sky130_fd_sc_hd__a21oi_1
XFILLER_138_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07235_ _08303_/A VGND VGND VPWR VPWR _08124_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_164_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07166_ _07166_/A _07166_/B VGND VGND VPWR VPWR _07205_/A sky130_fd_sc_hd__xnor2_1
XFILLER_118_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06117_ _14200_/Q _14198_/Q _14209_/Q VGND VGND VPWR VPWR _06117_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07097_ _07067_/A _07069_/B _07067_/B VGND VGND VPWR VPWR _07098_/B sky130_fd_sc_hd__o21ba_1
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06048_ _13975_/Q _13973_/Q _13977_/Q VGND VGND VPWR VPWR _06049_/B sky130_fd_sc_hd__mux2_1
XFILLER_160_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09807_ _09802_/B _09806_/Y _09834_/S VGND VGND VPWR VPWR _09808_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07999_ _13276_/Q _13277_/Q _13278_/Q _13279_/Q _08002_/B VGND VGND VPWR VPWR _07999_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_101_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09738_ _09673_/X _09732_/X _09734_/X _09737_/Y VGND VGND VPWR VPWR _09739_/B sky130_fd_sc_hd__o211a_1
XFILLER_27_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _13701_/Q VGND VGND VPWR VPWR _09883_/B sky130_fd_sc_hd__buf_4
XFILLER_15_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _14032_/Q _11510_/X _11700_/S VGND VGND VPWR VPWR _11701_/A sky130_fd_sc_hd__mux2_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _13799_/CLK _12680_/D VGND VGND VPWR VPWR _12680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11631_ _11631_/A VGND VGND VPWR VPWR _13991_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11562_ _11562_/A VGND VGND VPWR VPWR _13863_/D sky130_fd_sc_hd__clkbuf_1
X_14350_ _14697_/CLK hold16/X VGND VGND VPWR VPWR hold474/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10513_ _10511_/Y _10521_/B _10519_/A VGND VGND VPWR VPWR _10514_/A sky130_fd_sc_hd__mux2_1
X_13301_ _13303_/CLK hold111/X VGND VGND VPWR VPWR _13301_/Q sky130_fd_sc_hd__dfxtp_1
X_14281_ _14292_/CLK hold264/X VGND VGND VPWR VPWR _14281_/Q sky130_fd_sc_hd__dfxtp_1
X_11493_ _11493_/A VGND VGND VPWR VPWR _13832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13232_ _13617_/CLK hold57/X VGND VGND VPWR VPWR _13232_/Q sky130_fd_sc_hd__dfxtp_1
X_10444_ hold186/A _10444_/B _10449_/A VGND VGND VPWR VPWR _10453_/A sky130_fd_sc_hd__and3_1
XFILLER_108_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13163_ _13423_/CLK _13163_/D repeater57/X VGND VGND VPWR VPWR _13163_/Q sky130_fd_sc_hd__dfrtp_1
X_10375_ _10432_/A _10423_/A _10413_/B _10432_/B VGND VGND VPWR VPWR _10377_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_3_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12114_ _12114_/A VGND VGND VPWR VPWR _14472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13094_ _13587_/CLK hold297/X VGND VGND VPWR VPWR _13094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12045_ _12045_/A VGND VGND VPWR VPWR _14441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13996_ _14721_/CLK _13996_/D VGND VGND VPWR VPWR _13996_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12947_ _13280_/CLK _12947_/D VGND VGND VPWR VPWR hold318/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _12885_/CLK _12878_/D hold1/X VGND VGND VPWR VPWR _12878_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ _14617_/CLK _14617_/D VGND VGND VPWR VPWR _14617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11829_ _11829_/A VGND VGND VPWR VPWR _14106_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14548_ _14721_/CLK _14548_/D VGND VGND VPWR VPWR _14548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14479_ _14543_/CLK _14479_/D VGND VGND VPWR VPWR _14479_/Q sky130_fd_sc_hd__dfxtp_1
X_07020_ _13036_/D _07020_/B VGND VGND VPWR VPWR _07020_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_134_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08971_ _08971_/A _08971_/B VGND VGND VPWR VPWR _08972_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07922_ _13268_/Q _07947_/B VGND VGND VPWR VPWR _07923_/B sky130_fd_sc_hd__or2_1
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_69_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07853_ _13260_/Q _07853_/B _07853_/C VGND VGND VPWR VPWR _07885_/A sky130_fd_sc_hd__and3_1
XFILLER_84_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06804_ _06794_/B _06826_/B _06826_/A VGND VGND VPWR VPWR _06806_/B sky130_fd_sc_hd__a21o_1
XFILLER_110_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07784_ _07760_/A _07787_/C _07779_/A VGND VGND VPWR VPWR _07790_/A sky130_fd_sc_hd__a21o_1
XFILLER_72_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09523_ _09513_/A _09514_/X _09519_/B VGND VGND VPWR VPWR _09523_/X sky130_fd_sc_hd__a21bo_1
X_06735_ _06630_/A _06852_/B _06668_/X _06672_/X _06783_/S _06745_/A VGND VGND VPWR
+ VPWR _06736_/B sky130_fd_sc_hd__mux4_1
XFILLER_24_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09454_ _09454_/A _09454_/B _09454_/C _09454_/D VGND VGND VPWR VPWR _09455_/C sky130_fd_sc_hd__or4_1
X_06666_ _06659_/B _06661_/B _06659_/A VGND VGND VPWR VPWR _06681_/A sky130_fd_sc_hd__o21ba_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08405_ _08405_/A VGND VGND VPWR VPWR _12734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09385_ _09385_/A _09385_/B VGND VGND VPWR VPWR _09385_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_52_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06597_ _06597_/A _06597_/B VGND VGND VPWR VPWR _12898_/D sky130_fd_sc_hd__nor2_1
XFILLER_33_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08336_ _13382_/Q _13383_/Q VGND VGND VPWR VPWR _08340_/D sky130_fd_sc_hd__and2_1
XFILLER_137_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08267_ _08267_/A _08267_/B VGND VGND VPWR VPWR _08267_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_140_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _14153_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07218_ _07215_/Y _13036_/D _07218_/S VGND VGND VPWR VPWR _07219_/A sky130_fd_sc_hd__mux2_1
X_08198_ _08261_/A _10306_/A _13477_/Q _08177_/A VGND VGND VPWR VPWR _08199_/C sky130_fd_sc_hd__a31o_1
XFILLER_118_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07149_ _07149_/A _07175_/B VGND VGND VPWR VPWR _07150_/B sky130_fd_sc_hd__xnor2_2
XFILLER_118_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10160_ _10103_/A _14286_/D _10159_/X VGND VGND VPWR VPWR _10160_/X sky130_fd_sc_hd__a21o_1
XFILLER_105_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10091_ _10091_/A VGND VGND VPWR VPWR _13905_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13850_ _14180_/CLK _13850_/D VGND VGND VPWR VPWR _13850_/Q sky130_fd_sc_hd__dfxtp_1
X_12801_ _14275_/CLK _12801_/D VGND VGND VPWR VPWR hold438/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10993_ _10993_/A VGND VGND VPWR VPWR _10993_/X sky130_fd_sc_hd__clkbuf_4
X_13781_ _14647_/CLK _13781_/D VGND VGND VPWR VPWR _13781_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _13617_/CLK _12732_/D VGND VGND VPWR VPWR hold362/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _14702_/CLK _12663_/D VGND VGND VPWR VPWR _13244_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_31_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _14410_/CLK _14402_/D VGND VGND VPWR VPWR _14402_/Q sky130_fd_sc_hd__dfxtp_1
X_11614_ _11636_/A VGND VGND VPWR VPWR _11623_/S sky130_fd_sc_hd__buf_2
X_12594_ _12592_/X _12633_/B VGND VGND VPWR VPWR _12595_/A sky130_fd_sc_hd__and2b_1
XFILLER_11_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14333_ _14333_/CLK hold15/X VGND VGND VPWR VPWR hold221/A sky130_fd_sc_hd__dfxtp_1
X_11545_ _11545_/A VGND VGND VPWR VPWR _13855_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_131_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _14179_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11476_ _13827_/Q _11475_/X _11479_/S VGND VGND VPWR VPWR _11477_/A sky130_fd_sc_hd__mux2_1
X_14264_ _14656_/CLK _14264_/D VGND VGND VPWR VPWR _14264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10427_ _10431_/B _10427_/B VGND VGND VPWR VPWR _10428_/A sky130_fd_sc_hd__and2_1
X_13215_ _13366_/CLK hold493/X VGND VGND VPWR VPWR _13215_/Q sky130_fd_sc_hd__dfxtp_1
X_14195_ _14196_/CLK _14195_/D VGND VGND VPWR VPWR _14195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13146_ _13535_/CLK _13146_/D _12609_/A VGND VGND VPWR VPWR _13146_/Q sky130_fd_sc_hd__dfrtp_1
X_10358_ _10358_/A VGND VGND VPWR VPWR _12987_/D sky130_fd_sc_hd__clkbuf_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _13528_/CLK hold294/X VGND VGND VPWR VPWR _13077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10289_ hold500/A VGND VGND VPWR VPWR hold506/A sky130_fd_sc_hd__clkinv_2
X_12028_ _14681_/Q _12034_/B _12030_/C VGND VGND VPWR VPWR _12029_/A sky130_fd_sc_hd__and3_1
XFILLER_78_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13979_ _14533_/CLK _13979_/D VGND VGND VPWR VPWR _13979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06520_ _06520_/A _06520_/B VGND VGND VPWR VPWR _06520_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_80_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06451_ _06436_/A _06433_/A _06436_/B _06450_/X VGND VGND VPWR VPWR _06452_/B sky130_fd_sc_hd__a31oi_4
XFILLER_22_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09170_ _09177_/A _09177_/B VGND VGND VPWR VPWR _09172_/A sky130_fd_sc_hd__nor2_1
X_06382_ _14431_/Q hold187/A _06425_/S VGND VGND VPWR VPWR _06382_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08121_ _08199_/A _08120_/C _13355_/Q VGND VGND VPWR VPWR _08121_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_122_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _13626_/CLK sky130_fd_sc_hd__clkbuf_16
X_08052_ _08052_/A VGND VGND VPWR VPWR _12687_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07003_ _13029_/Q _08020_/B VGND VGND VPWR VPWR _07003_/Y sky130_fd_sc_hd__nand2_1
XFILLER_134_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08954_ _08954_/A _08954_/B VGND VGND VPWR VPWR _08993_/A sky130_fd_sc_hd__xnor2_1
XFILLER_88_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07905_ _07905_/A _07905_/B VGND VGND VPWR VPWR _07906_/B sky130_fd_sc_hd__nor2_1
X_08885_ _08855_/A _08857_/B _08855_/B VGND VGND VPWR VPWR _08886_/B sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_189_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _14726_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07836_ _07835_/A _07858_/A _07858_/B VGND VGND VPWR VPWR _07836_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07767_ _07738_/Y _07766_/X _07781_/S VGND VGND VPWR VPWR _07768_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09506_ _09506_/A VGND VGND VPWR VPWR _09506_/X sky130_fd_sc_hd__clkbuf_2
X_06718_ _06719_/A _06716_/Y _06720_/C _06881_/A VGND VGND VPWR VPWR _06733_/B sky130_fd_sc_hd__a22o_1
X_07698_ _13114_/Q VGND VGND VPWR VPWR _07772_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09437_ _09502_/A VGND VGND VPWR VPWR _09437_/X sky130_fd_sc_hd__clkbuf_2
X_06649_ _13038_/Q VGND VGND VPWR VPWR _06674_/C sky130_fd_sc_hd__buf_2
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09368_ _09367_/B _09367_/C _13590_/Q VGND VGND VPWR VPWR _09368_/X sky130_fd_sc_hd__a21o_1
X_08319_ _08325_/D _08319_/B VGND VGND VPWR VPWR _13377_/D sky130_fd_sc_hd__nor2_1
XFILLER_21_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_113_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _13377_/CLK sky130_fd_sc_hd__clkbuf_16
X_09299_ _13288_/Q _13526_/Q _09299_/S VGND VGND VPWR VPWR _09300_/A sky130_fd_sc_hd__mux2_1
XANTENNA_60 input8/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_71 _13552_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11330_ _11330_/A VGND VGND VPWR VPWR _11355_/S sky130_fd_sc_hd__buf_2
XANTENNA_82 _11636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 _13544_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11261_ _14280_/Q _14671_/Q _13778_/Q _14726_/Q _10914_/A _10918_/A VGND VGND VPWR
+ VPWR _11262_/B sky130_fd_sc_hd__mux4_1
X_10212_ _14095_/Q _14079_/Q _14384_/D VGND VGND VPWR VPWR _10213_/A sky130_fd_sc_hd__mux2_1
X_13000_ _13525_/CLK _13000_/D hold1/X VGND VGND VPWR VPWR _13000_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11192_ _11240_/A _11192_/B VGND VGND VPWR VPWR _11192_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10143_ _10143_/A VGND VGND VPWR VPWR _10143_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10074_ _14044_/D _10073_/X _14049_/D VGND VGND VPWR VPWR _10074_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13902_ _14050_/CLK _13902_/D VGND VGND VPWR VPWR hold286/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13833_ _14707_/CLK _13833_/D VGND VGND VPWR VPWR _13833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13764_ _14712_/CLK _13764_/D VGND VGND VPWR VPWR _13764_/Q sky130_fd_sc_hd__dfxtp_1
X_10976_ _11035_/A _10976_/B VGND VGND VPWR VPWR _10976_/Y sky130_fd_sc_hd__nor2_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12715_ _13596_/CLK _12715_/D VGND VGND VPWR VPWR hold483/A sky130_fd_sc_hd__dfxtp_1
X_13695_ _13855_/CLK _13695_/D repeater57/X VGND VGND VPWR VPWR _13695_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_70_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12646_ _14742_/Q _12567_/X _12645_/X _12609_/X VGND VGND VPWR VPWR _14747_/D sky130_fd_sc_hd__o211a_1
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_104_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _13602_/CLK sky130_fd_sc_hd__clkbuf_16
X_12577_ _12573_/Y _11655_/A _11712_/B _12625_/A _12576_/X VGND VGND VPWR VPWR _12577_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_12_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14316_ _14617_/CLK _14316_/D VGND VGND VPWR VPWR _14316_/Q sky130_fd_sc_hd__dfxtp_1
X_11528_ _11528_/A VGND VGND VPWR VPWR _13848_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold308 hold308/A VGND VGND VPWR VPWR hold308/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold319 hold319/A VGND VGND VPWR VPWR hold319/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14247_ _14250_/CLK _14247_/D VGND VGND VPWR VPWR _14247_/Q sky130_fd_sc_hd__dfxtp_1
X_11459_ _14697_/Q VGND VGND VPWR VPWR _11459_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14178_ _14196_/CLK _14178_/D VGND VGND VPWR VPWR _14178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _13434_/CLK hold59/X VGND VGND VPWR VPWR hold210/A sky130_fd_sc_hd__dfxtp_1
XFILLER_140_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05951_ _13864_/Q _13865_/Q _05951_/C _05951_/D VGND VGND VPWR VPWR _05952_/B sky130_fd_sc_hd__and4_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08670_ _08629_/X _08641_/A _08653_/B _08664_/C _08669_/X VGND VGND VPWR VPWR _08689_/B
+ sky130_fd_sc_hd__o41ai_4
XFILLER_54_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07621_ _13246_/D VGND VGND VPWR VPWR _07747_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07552_ _07553_/B _07553_/C _07559_/A VGND VGND VPWR VPWR _07556_/B sky130_fd_sc_hd__a21o_1
XFILLER_53_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06503_ _10346_/A _13109_/D VGND VGND VPWR VPWR _06554_/C sky130_fd_sc_hd__nor2_2
XFILLER_22_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07483_ _07493_/A _07483_/B VGND VGND VPWR VPWR _07504_/B sky130_fd_sc_hd__nand2_1
XFILLER_61_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09222_ _09195_/A _09242_/B _09244_/A VGND VGND VPWR VPWR _09223_/B sky130_fd_sc_hd__o21ba_1
X_06434_ _06482_/A _06513_/B _06417_/X _06471_/A _12878_/Q VGND VGND VPWR VPWR _06434_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_139_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09153_ _13534_/Q _09153_/B _09153_/C VGND VGND VPWR VPWR _09159_/C sky130_fd_sc_hd__and3_1
X_06365_ _14645_/Q _14428_/D VGND VGND VPWR VPWR _06365_/Y sky130_fd_sc_hd__nor2_1
X_08104_ _08162_/B VGND VGND VPWR VPWR _08208_/A sky130_fd_sc_hd__inv_2
XFILLER_108_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09084_ _09084_/A _13523_/Q VGND VGND VPWR VPWR _09085_/B sky130_fd_sc_hd__nand2_1
X_06296_ _14162_/Q _14206_/D VGND VGND VPWR VPWR _06296_/X sky130_fd_sc_hd__and2_1
XFILLER_147_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08035_ _08035_/A VGND VGND VPWR VPWR _12676_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09986_ _09986_/A VGND VGND VPWR VPWR _13706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08937_ _08937_/A _08963_/B VGND VGND VPWR VPWR _08938_/B sky130_fd_sc_hd__xnor2_1
XFILLER_69_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08868_ _08843_/Y _08867_/Y _11268_/A VGND VGND VPWR VPWR _08869_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07819_ _13255_/Q _07819_/B VGND VGND VPWR VPWR _07820_/B sky130_fd_sc_hd__and2_1
XFILLER_29_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08799_ _13515_/D VGND VGND VPWR VPWR _08819_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_44_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10830_ _10830_/A VGND VGND VPWR VPWR _13176_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10761_ _10761_/A VGND VGND VPWR VPWR _13044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12500_ _12502_/A _12502_/B hold464/X VGND VGND VPWR VPWR _12501_/A sky130_fd_sc_hd__and3_1
XFILLER_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10692_ _12882_/Q _10698_/B VGND VGND VPWR VPWR _10693_/A sky130_fd_sc_hd__and2_1
X_13480_ _14251_/CLK hold185/X VGND VGND VPWR VPWR _13480_/Q sky130_fd_sc_hd__dfxtp_1
X_12431_ _14648_/Q _14694_/Q _12439_/S VGND VGND VPWR VPWR _12432_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12362_ _14604_/Q _11978_/X _12364_/S VGND VGND VPWR VPWR _12363_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14101_ _14319_/CLK _14101_/D VGND VGND VPWR VPWR _14101_/Q sky130_fd_sc_hd__dfxtp_1
X_11313_ _14515_/Q VGND VGND VPWR VPWR _11313_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_153_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12293_ _12315_/A VGND VGND VPWR VPWR _12302_/S sky130_fd_sc_hd__buf_2
XFILLER_154_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11244_ _14317_/Q _14487_/Q _14243_/Q _14073_/Q _11208_/X _11209_/X VGND VGND VPWR
+ VPWR _11244_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14032_ _14722_/CLK _14032_/D VGND VGND VPWR VPWR _14032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11175_ _11175_/A VGND VGND VPWR VPWR _11175_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10126_ _10126_/A VGND VGND VPWR VPWR _14177_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10057_ _13920_/Q _10056_/X _10060_/A VGND VGND VPWR VPWR _10057_/X sky130_fd_sc_hd__a21o_1
XFILLER_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13816_ _14633_/CLK _13816_/D VGND VGND VPWR VPWR hold324/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13747_ _14588_/CLK _13747_/D VGND VGND VPWR VPWR _13747_/Q sky130_fd_sc_hd__dfxtp_2
X_10959_ _14258_/Q _14649_/Q _13756_/Q _14704_/Q _10940_/X _10942_/X VGND VGND VPWR
+ VPWR _10960_/B sky130_fd_sc_hd__mux4_1
X_13678_ _13680_/CLK _13678_/D repeater56/X VGND VGND VPWR VPWR _13678_/Q sky130_fd_sc_hd__dfrtp_1
X_12629_ _12631_/B _12631_/C _12641_/A VGND VGND VPWR VPWR _12629_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06150_ _06289_/S VGND VGND VPWR VPWR _10110_/A sky130_fd_sc_hd__clkbuf_2
X_06081_ _13946_/Q _13938_/Q _10023_/A VGND VGND VPWR VPWR _10606_/A sky130_fd_sc_hd__mux2_1
Xhold105 hold105/A VGND VGND VPWR VPWR hold105/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold116 hold116/A VGND VGND VPWR VPWR hold116/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold127 hold127/A VGND VGND VPWR VPWR hold127/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold138 hold138/A VGND VGND VPWR VPWR hold138/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold149 hold149/A VGND VGND VPWR VPWR hold149/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ _09840_/A VGND VGND VPWR VPWR _09840_/Y sky130_fd_sc_hd__inv_2
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _09749_/A _09761_/A _09761_/B VGND VGND VPWR VPWR _09771_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_140_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06983_ _06968_/A _06968_/B _06981_/Y _06982_/X VGND VGND VPWR VPWR _06996_/A sky130_fd_sc_hd__a31oi_2
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08722_ _09524_/B VGND VGND VPWR VPWR _09530_/B sky130_fd_sc_hd__buf_2
X_05934_ _05934_/A _05934_/B _05934_/C VGND VGND VPWR VPWR _05935_/C sky130_fd_sc_hd__or3_1
XFILLER_39_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08653_ _08653_/A _08653_/B VGND VGND VPWR VPWR _08654_/B sky130_fd_sc_hd__or2_1
XFILLER_81_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07604_ _07800_/S VGND VGND VPWR VPWR _11266_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08584_ _08567_/A _08582_/B _08567_/C _08581_/B VGND VGND VPWR VPWR _09424_/C sky130_fd_sc_hd__a31o_1
XFILLER_54_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07535_ _07477_/B _07533_/Y _07534_/X _07507_/X VGND VGND VPWR VPWR _07548_/A sky130_fd_sc_hd__a211o_2
XFILLER_23_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07466_ _09207_/B VGND VGND VPWR VPWR _09212_/B sky130_fd_sc_hd__buf_2
XFILLER_139_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09205_ _09205_/A _09201_/B VGND VGND VPWR VPWR _09210_/B sky130_fd_sc_hd__or2b_1
X_06417_ _06427_/S _06415_/X _06416_/X _10346_/A VGND VGND VPWR VPWR _06417_/X sky130_fd_sc_hd__a211o_1
X_07397_ _07343_/X _07394_/X _07396_/X VGND VGND VPWR VPWR _13141_/D sky130_fd_sc_hd__a21o_1
X_06348_ _14406_/D _14407_/D _14408_/D _06348_/D VGND VGND VPWR VPWR _06348_/X sky130_fd_sc_hd__and4_1
X_09136_ _09161_/A _09137_/B _07524_/X VGND VGND VPWR VPWR _09136_/X sky130_fd_sc_hd__a21o_1
XFILLER_148_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09067_ _13231_/Q _13460_/Q _09075_/S VGND VGND VPWR VPWR _09068_/A sky130_fd_sc_hd__mux2_1
X_06279_ _13812_/Q _13796_/Q _06281_/S VGND VGND VPWR VPWR _06280_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08018_ _08018_/A _08018_/B _08018_/C VGND VGND VPWR VPWR _08018_/Y sky130_fd_sc_hd__nand3_1
XFILLER_2_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09969_ _09969_/A VGND VGND VPWR VPWR _12870_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12980_ _13280_/CLK hold318/X VGND VGND VPWR VPWR _12980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11931_ _11931_/A VGND VGND VPWR VPWR _11940_/S sky130_fd_sc_hd__buf_2
XFILLER_57_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _14705_/CLK _14650_/D VGND VGND VPWR VPWR _14650_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _14229_/Q _11475_/X _11864_/S VGND VGND VPWR VPWR _11863_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _13621_/CLK _13601_/D repeater56/X VGND VGND VPWR VPWR _13601_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10813_ _10813_/A VGND VGND VPWR VPWR _13068_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _14619_/CLK _14581_/D VGND VGND VPWR VPWR _14581_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11793_ _13568_/Q _11795_/B VGND VGND VPWR VPWR _11794_/A sky130_fd_sc_hd__and2_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13532_ _13532_/CLK _13532_/D repeater57/X VGND VGND VPWR VPWR _13532_/Q sky130_fd_sc_hd__dfrtp_2
X_10744_ _12906_/Q _10748_/B VGND VGND VPWR VPWR _10745_/A sky130_fd_sc_hd__and2_1
XFILLER_13_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13463_ _13622_/CLK _13463_/D repeater57/X VGND VGND VPWR VPWR _13463_/Q sky130_fd_sc_hd__dfrtp_1
X_10675_ _14343_/Q _10671_/X _10656_/X VGND VGND VPWR VPWR _10675_/Y sky130_fd_sc_hd__a21boi_1
X_12414_ _12418_/A _12418_/B input2/X VGND VGND VPWR VPWR _12415_/A sky130_fd_sc_hd__and3_1
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13394_ _13593_/CLK hold458/X VGND VGND VPWR VPWR _13394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12345_ _14596_/Q _11950_/X _12353_/S VGND VGND VPWR VPWR _12346_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12276_ _11370_/X _14553_/Q _12278_/S VGND VGND VPWR VPWR _12277_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14015_ _14533_/CLK _14015_/D VGND VGND VPWR VPWR _14015_/Q sky130_fd_sc_hd__dfxtp_1
X_11227_ _11227_/A VGND VGND VPWR VPWR _11227_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11158_ _11136_/X _11151_/X _11156_/X _11157_/X VGND VGND VPWR VPWR _11158_/X sky130_fd_sc_hd__o211a_1
XFILLER_122_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10109_ _14180_/Q _14172_/Q _10110_/A VGND VGND VPWR VPWR _10616_/C sky130_fd_sc_hd__mux2_1
X_11089_ _14606_/Q _14568_/Q _14499_/Q _14451_/Q _11044_/X _11045_/X VGND VGND VPWR
+ VPWR _11090_/A sky130_fd_sc_hd__mux4_1
XFILLER_49_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07320_ _07320_/A VGND VGND VPWR VPWR _07321_/A sky130_fd_sc_hd__inv_2
XFILLER_32_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07251_ _07311_/A VGND VGND VPWR VPWR _07461_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06202_ _06202_/A VGND VGND VPWR VPWR _14368_/D sky130_fd_sc_hd__clkbuf_1
X_07182_ _07182_/A _07182_/B _07182_/C VGND VGND VPWR VPWR _07183_/B sky130_fd_sc_hd__and3_1
X_06133_ _14205_/Q _14203_/Q _10107_/A VGND VGND VPWR VPWR _06133_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06064_ _06063_/X _06060_/X _10019_/A VGND VGND VPWR VPWR _06065_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09823_ _09815_/A _09816_/A _09815_/B _09812_/A VGND VGND VPWR VPWR _09824_/B sky130_fd_sc_hd__a31o_1
XFILLER_101_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09754_ _09748_/B _09753_/X _09774_/S VGND VGND VPWR VPWR _09755_/A sky130_fd_sc_hd__mux2_1
X_06966_ _13022_/Q _13023_/Q _06895_/B VGND VGND VPWR VPWR _06973_/B sky130_fd_sc_hd__o21ai_1
XFILLER_74_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08705_ _08617_/X _08709_/B _08704_/Y _08696_/X VGND VGND VPWR VPWR _13453_/D sky130_fd_sc_hd__a31o_1
X_05917_ _13734_/Q _13735_/Q _13736_/Q _05917_/D VGND VGND VPWR VPWR _05917_/X sky130_fd_sc_hd__and4_1
X_09685_ _14218_/Q _14216_/Q _09688_/S VGND VGND VPWR VPWR _09685_/X sky130_fd_sc_hd__mux2_1
X_06897_ _07932_/A VGND VGND VPWR VPWR _06897_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _13702_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08636_ _08546_/Y _08635_/Y _08544_/X VGND VGND VPWR VPWR _09457_/C sky130_fd_sc_hd__o21ai_4
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ _08567_/A _08582_/B _08567_/C VGND VGND VPWR VPWR _09414_/B sky130_fd_sc_hd__nand3_1
XFILLER_42_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07518_ _07495_/X _07516_/X _07517_/Y _07499_/X VGND VGND VPWR VPWR _13152_/D sky130_fd_sc_hd__a31o_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08498_ _08512_/A _08497_/Y VGND VGND VPWR VPWR _08500_/A sky130_fd_sc_hd__or2b_1
XFILLER_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07449_ _13146_/Q _07450_/A VGND VGND VPWR VPWR _07452_/A sky130_fd_sc_hd__and2_1
X_10460_ _10460_/A _10485_/A VGND VGND VPWR VPWR _10462_/A sky130_fd_sc_hd__nand2_1
XFILLER_164_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09119_ _13528_/Q _09120_/B VGND VGND VPWR VPWR _09119_/Y sky130_fd_sc_hd__nand2_1
X_10391_ _10407_/A _10391_/B VGND VGND VPWR VPWR _10393_/B sky130_fd_sc_hd__nor2_1
X_12130_ _12130_/A VGND VGND VPWR VPWR _12139_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_108_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12061_ _11307_/X _14449_/Q _12063_/S VGND VGND VPWR VPWR _12062_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold480 data_i[1] VGND VGND VPWR VPWR input12/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold491 hold10/X VGND VGND VPWR VPWR hold491/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11012_ _14018_/Q _13984_/Q _13824_/Q _14536_/Q _11010_/X _11011_/X VGND VGND VPWR
+ VPWR _11014_/A sky130_fd_sc_hd__mux4_1
XFILLER_104_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12963_ _13263_/CLK hold112/X VGND VGND VPWR VPWR _12963_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_84_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _14010_/CLK sky130_fd_sc_hd__clkbuf_16
X_14702_ _14702_/CLK _14702_/D VGND VGND VPWR VPWR _14702_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11914_ _14264_/Q _11472_/X _11918_/S VGND VGND VPWR VPWR _11915_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _12970_/CLK _12894_/D hold1/X VGND VGND VPWR VPWR _12894_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _14633_/CLK _14633_/D VGND VGND VPWR VPWR _14633_/Q sky130_fd_sc_hd__dfxtp_1
X_11845_ _14221_/Q _11446_/X _11853_/S VGND VGND VPWR VPWR _11846_/A sky130_fd_sc_hd__mux2_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _14602_/CLK _14564_/D VGND VGND VPWR VPWR _14564_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11776_ _13560_/Q _11784_/B VGND VGND VPWR VPWR _11777_/A sky130_fd_sc_hd__and2_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13515_ _13520_/CLK _13515_/D VGND VGND VPWR VPWR _14211_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_14_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10727_ _12898_/Q _10731_/B VGND VGND VPWR VPWR _10728_/A sky130_fd_sc_hd__and2_1
XFILLER_159_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14495_ _14495_/CLK _14495_/D VGND VGND VPWR VPWR _14495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13446_ _13598_/CLK _13446_/D repeater56/X VGND VGND VPWR VPWR _13446_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_127_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10658_ _14337_/Q _14334_/Q _10657_/Y VGND VGND VPWR VPWR _12912_/D sky130_fd_sc_hd__a21oi_2
XFILLER_155_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13377_ _13377_/CLK _13377_/D _12609_/A VGND VGND VPWR VPWR _13377_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10589_ _13467_/Q _13472_/Q _13470_/Q _08464_/X VGND VGND VPWR VPWR _13467_/D sky130_fd_sc_hd__o31a_1
X_12328_ _14579_/Q _12019_/X _12332_/S VGND VGND VPWR VPWR _12329_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12259_ _11326_/X _14545_/Q _12259_/S VGND VGND VPWR VPWR _12260_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06820_ _06820_/A _06820_/B _06820_/C VGND VGND VPWR VPWR _06820_/Y sky130_fd_sc_hd__nand3_1
XFILLER_96_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06751_ _06782_/A _06751_/B VGND VGND VPWR VPWR _06751_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_75_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _14012_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_48_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09470_ _09475_/B _09469_/Y _08655_/X VGND VGND VPWR VPWR _13603_/D sky130_fd_sc_hd__a21o_1
X_06682_ _06681_/B _06681_/C _06681_/A VGND VGND VPWR VPWR _06682_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08421_ _13105_/Q _13386_/Q _09299_/S VGND VGND VPWR VPWR _08422_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08352_ _13468_/D VGND VGND VPWR VPWR _08397_/A sky130_fd_sc_hd__clkbuf_4
X_07303_ _13135_/Q _09113_/B VGND VGND VPWR VPWR _07305_/B sky130_fd_sc_hd__xnor2_1
XFILLER_32_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08283_ _08283_/A VGND VGND VPWR VPWR _08283_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07234_ _13165_/Q VGND VGND VPWR VPWR _08303_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07165_ _07165_/A _07190_/D VGND VGND VPWR VPWR _07166_/B sky130_fd_sc_hd__nand2_1
XFILLER_106_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06116_ _14201_/Q _14199_/Q _14209_/Q VGND VGND VPWR VPWR _06116_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07096_ _07126_/A _07126_/B VGND VGND VPWR VPWR _07098_/A sky130_fd_sc_hd__xnor2_1
XFILLER_161_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06047_ _13968_/Q _13966_/Q _13977_/Q VGND VGND VPWR VPWR _06047_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09806_ _09806_/A _09806_/B VGND VGND VPWR VPWR _09806_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07998_ _07998_/A _07998_/B VGND VGND VPWR VPWR _07998_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09737_ _09836_/A _09778_/A _09675_/X _13703_/Q VGND VGND VPWR VPWR _09737_/Y sky130_fd_sc_hd__a31oi_1
X_06949_ _06945_/X _06947_/Y _06948_/X _06907_/X VGND VGND VPWR VPWR _13021_/D sky130_fd_sc_hd__a31o_1
XFILLER_28_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_66_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _13359_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09668_ _09778_/B _09678_/C VGND VGND VPWR VPWR _09671_/A sky130_fd_sc_hd__nand2_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _08620_/C _08618_/X VGND VGND VPWR VPWR _08630_/B sky130_fd_sc_hd__or2b_1
XFILLER_131_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _09599_/A VGND VGND VPWR VPWR _12814_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _13991_/Q _11488_/X _11634_/S VGND VGND VPWR VPWR _11631_/A sky130_fd_sc_hd__mux2_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11561_ _13639_/Q _11563_/B VGND VGND VPWR VPWR _11562_/A sky130_fd_sc_hd__and2_1
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13300_ _13303_/CLK hold418/X VGND VGND VPWR VPWR _13300_/Q sky130_fd_sc_hd__dfxtp_1
X_10512_ _10512_/A _12991_/D VGND VGND VPWR VPWR _10519_/A sky130_fd_sc_hd__and2_1
XFILLER_128_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14280_ _14725_/CLK _14280_/D VGND VGND VPWR VPWR _14280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11492_ _13832_/Q _11491_/X _11495_/S VGND VGND VPWR VPWR _11493_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13231_ _13617_/CLK hold447/X VGND VGND VPWR VPWR _13231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10443_ _10443_/A VGND VGND VPWR VPWR _14006_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13162_ _13554_/CLK _13162_/D _12609_/A VGND VGND VPWR VPWR _13162_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10374_ _10374_/A VGND VGND VPWR VPWR _10413_/B sky130_fd_sc_hd__inv_2
XFILLER_151_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12113_ _14472_/Q _11975_/X _12117_/S VGND VGND VPWR VPWR _12114_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13093_ _13587_/CLK hold404/X VGND VGND VPWR VPWR _13093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12044_ _11272_/X _14441_/Q _12052_/S VGND VGND VPWR VPWR _12045_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13995_ _14720_/CLK _13995_/D VGND VGND VPWR VPWR _13995_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_57_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _14634_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_58_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ _13280_/CLK _12946_/D VGND VGND VPWR VPWR hold285/A sky130_fd_sc_hd__dfxtp_1
XFILLER_65_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ _12885_/CLK _12877_/D hold1/X VGND VGND VPWR VPWR _12877_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _14617_/CLK _14616_/D VGND VGND VPWR VPWR _14616_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _13584_/Q _11828_/B VGND VGND VPWR VPWR _11829_/A sky130_fd_sc_hd__and2_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _14720_/CLK _14547_/D VGND VGND VPWR VPWR _14547_/Q sky130_fd_sc_hd__dfxtp_1
X_11759_ _11759_/A VGND VGND VPWR VPWR _14070_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14478_ _14652_/CLK _14478_/D VGND VGND VPWR VPWR _14478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13429_ _14588_/CLK hold71/X VGND VGND VPWR VPWR _13429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08970_ _08970_/A _08970_/B _08970_/C VGND VGND VPWR VPWR _08971_/B sky130_fd_sc_hd__and3_1
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07921_ _13268_/Q _07955_/B VGND VGND VPWR VPWR _07923_/A sky130_fd_sc_hd__nand2_1
X_07852_ _07852_/A VGND VGND VPWR VPWR _13259_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06803_ _13006_/Q _06781_/B _06791_/A VGND VGND VPWR VPWR _06826_/B sky130_fd_sc_hd__a21oi_1
Xinput1 data_i[0] VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_6
X_07783_ _07783_/A VGND VGND VPWR VPWR _07787_/C sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_48_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _14680_/CLK sky130_fd_sc_hd__clkbuf_16
X_09522_ _09520_/Y _09521_/X _08735_/X VGND VGND VPWR VPWR _13610_/D sky130_fd_sc_hd__o21bai_1
X_06734_ _06703_/X _06731_/Y _06733_/X VGND VGND VPWR VPWR _13003_/D sky130_fd_sc_hd__o21bai_1
XFILLER_24_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09453_ _09455_/B _09446_/X _09449_/Y _09455_/A VGND VGND VPWR VPWR _09460_/B sky130_fd_sc_hd__a31o_1
X_06665_ _07802_/A VGND VGND VPWR VPWR _06665_/X sky130_fd_sc_hd__buf_2
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08404_ _13098_/Q _13379_/Q _08406_/S VGND VGND VPWR VPWR _08405_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09384_ _09377_/A _09377_/B _09383_/X VGND VGND VPWR VPWR _09385_/B sky130_fd_sc_hd__a21o_1
XFILLER_51_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06596_ _12898_/Q _06593_/A _06542_/X VGND VGND VPWR VPWR _06597_/B sky130_fd_sc_hd__o21ai_1
X_08335_ _13382_/Q _08333_/A _08334_/Y VGND VGND VPWR VPWR _13382_/D sky130_fd_sc_hd__a21oi_1
XFILLER_138_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08266_ _08256_/A _08257_/A _08256_/B _08253_/A VGND VGND VPWR VPWR _08267_/B sky130_fd_sc_hd__a31o_1
X_07217_ _07217_/A VGND VGND VPWR VPWR _13352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08197_ _08197_/A VGND VGND VPWR VPWR _10306_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07148_ _07115_/A _07115_/B _07121_/A _07121_/B VGND VGND VPWR VPWR _07175_/B sky130_fd_sc_hd__a22o_1
XFILLER_106_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07079_ _07156_/A _07079_/B VGND VGND VPWR VPWR _07079_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10090_ _10086_/X _10089_/X _10095_/S VGND VGND VPWR VPWR _10091_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_39_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _13264_/CLK sky130_fd_sc_hd__clkbuf_16
X_12800_ _14275_/CLK _12800_/D VGND VGND VPWR VPWR hold375/A sky130_fd_sc_hd__dfxtp_1
XFILLER_90_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13780_ _14647_/CLK _13780_/D VGND VGND VPWR VPWR _13780_/Q sky130_fd_sc_hd__dfxtp_1
X_10992_ _11162_/A VGND VGND VPWR VPWR _10993_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _13617_/CLK _12731_/D VGND VGND VPWR VPWR hold492/A sky130_fd_sc_hd__dfxtp_1
XFILLER_83_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _14737_/CLK _12662_/D _12609_/A VGND VGND VPWR VPWR _12662_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _14410_/CLK _14401_/D VGND VGND VPWR VPWR _14401_/Q sky130_fd_sc_hd__dfxtp_1
X_11613_ _11613_/A VGND VGND VPWR VPWR _13983_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ _12609_/A VGND VGND VPWR VPWR _12633_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_129_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14332_ _14333_/CLK hold221/X VGND VGND VPWR VPWR hold78/A sky130_fd_sc_hd__dfxtp_1
XFILLER_128_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11544_ _13631_/Q _11552_/B VGND VGND VPWR VPWR _11545_/A sky130_fd_sc_hd__and2_1
XFILLER_7_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14263_ _14709_/CLK _14263_/D VGND VGND VPWR VPWR _14263_/Q sky130_fd_sc_hd__dfxtp_1
X_11475_ _14513_/Q VGND VGND VPWR VPWR _11475_/X sky130_fd_sc_hd__clkbuf_2
X_13214_ _13434_/CLK hold353/X VGND VGND VPWR VPWR _13214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10426_ _10426_/A _10426_/B _10426_/C VGND VGND VPWR VPWR _10427_/B sky130_fd_sc_hd__or3_1
XFILLER_136_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14194_ _14209_/CLK _14194_/D VGND VGND VPWR VPWR _14194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13145_ _13535_/CLK _13145_/D repeater57/X VGND VGND VPWR VPWR _13145_/Q sky130_fd_sc_hd__dfrtp_2
X_10357_ _10359_/B _10357_/B VGND VGND VPWR VPWR _10358_/A sky130_fd_sc_hd__or2_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13076_ _13076_/CLK _13076_/D VGND VGND VPWR VPWR _13076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10288_ hold49/A VGND VGND VPWR VPWR hold505/A sky130_fd_sc_hd__inv_2
XFILLER_39_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12027_ _12027_/A VGND VGND VPWR VPWR _14318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13978_ _13978_/CLK _13978_/D VGND VGND VPWR VPWR _13978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12929_ _13265_/CLK _12929_/D VGND VGND VPWR VPWR hold107/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06450_ _12879_/Q _06450_/B VGND VGND VPWR VPWR _06450_/X sky130_fd_sc_hd__and2_1
XFILLER_92_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06381_ _13106_/D VGND VGND VPWR VPWR _06425_/S sky130_fd_sc_hd__clkbuf_2
X_08120_ _08164_/A _13355_/Q _08120_/C VGND VGND VPWR VPWR _08122_/A sky130_fd_sc_hd__and3_1
X_08051_ _12963_/Q _13263_/Q _08051_/S VGND VGND VPWR VPWR _08052_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07002_ _06945_/X _07000_/X _07001_/Y _06974_/X VGND VGND VPWR VPWR _13028_/D sky130_fd_sc_hd__a31o_1
XFILLER_143_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08953_ _08953_/A _08978_/D VGND VGND VPWR VPWR _08954_/B sky130_fd_sc_hd__nand2_1
XFILLER_102_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07904_ _07904_/A _07904_/B VGND VGND VPWR VPWR _07905_/B sky130_fd_sc_hd__nor2_1
X_08884_ _08914_/A _08914_/B VGND VGND VPWR VPWR _08886_/A sky130_fd_sc_hd__xnor2_1
XFILLER_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07835_ _07835_/A _07858_/A _07858_/B VGND VGND VPWR VPWR _07835_/Y sky130_fd_sc_hd__nand3_1
XFILLER_56_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07766_ _07791_/A _07766_/B VGND VGND VPWR VPWR _07766_/X sky130_fd_sc_hd__xor2_1
XFILLER_71_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09505_ _09505_/A _09505_/B _09509_/D VGND VGND VPWR VPWR _09505_/Y sky130_fd_sc_hd__nand3_1
X_06717_ _06630_/A _06841_/B _06645_/X _06646_/X _06783_/S _06745_/A VGND VGND VPWR
+ VPWR _06720_/C sky130_fd_sc_hd__mux4_1
X_07697_ _07697_/A _07697_/B VGND VGND VPWR VPWR _07703_/A sky130_fd_sc_hd__xor2_1
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09436_ _08784_/X _09443_/B _09435_/Y _08603_/X VGND VGND VPWR VPWR _13599_/D sky130_fd_sc_hd__a31o_1
X_06648_ _06705_/S _12672_/Q VGND VGND VPWR VPWR _06648_/X sky130_fd_sc_hd__and2b_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09367_ _13590_/Q _09367_/B _09367_/C VGND VGND VPWR VPWR _09369_/A sky130_fd_sc_hd__and3_1
X_06579_ _06574_/X _06584_/D _06578_/Y _06586_/A VGND VGND VPWR VPWR _12893_/D sky130_fd_sc_hd__a211oi_1
X_08318_ _13377_/Q _08316_/A _08338_/A VGND VGND VPWR VPWR _08319_/B sky130_fd_sc_hd__o21ai_1
XANTENNA_50 hold499/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09298_ _09298_/A VGND VGND VPWR VPWR _12777_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_61 input8/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _13553_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 _12185_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08249_ _08249_/A VGND VGND VPWR VPWR _13365_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_94 input12/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11260_ _11260_/A VGND VGND VPWR VPWR _11260_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10211_ _06215_/D _06324_/Y _14414_/D _10203_/X VGND VGND VPWR VPWR _14422_/D sky130_fd_sc_hd__a22o_1
XFILLER_106_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11191_ _14274_/Q _14665_/Q _13772_/Q _14720_/Q _11162_/X _11163_/X VGND VGND VPWR
+ VPWR _11192_/B sky130_fd_sc_hd__mux4_1
XFILLER_122_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10142_ hold184/A _10143_/A _10147_/A VGND VGND VPWR VPWR _14283_/D sky130_fd_sc_hd__a21o_1
X_10073_ _10016_/A _14042_/D _10072_/X VGND VGND VPWR VPWR _10073_/X sky130_fd_sc_hd__a21o_1
XFILLER_153_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13901_ _14210_/CLK hold254/X VGND VGND VPWR VPWR hold225/A sky130_fd_sc_hd__dfxtp_1
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13832_ _14707_/CLK _13832_/D VGND VGND VPWR VPWR _13832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13763_ _14710_/CLK _13763_/D VGND VGND VPWR VPWR _13763_/Q sky130_fd_sc_hd__dfxtp_1
X_10975_ _14259_/Q _14650_/Q _13757_/Q _14705_/Q _10940_/X _10942_/X VGND VGND VPWR
+ VPWR _10976_/B sky130_fd_sc_hd__mux4_1
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12714_ _13596_/CLK _12714_/D VGND VGND VPWR VPWR hold475/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13694_ _13811_/CLK _13694_/D repeater57/X VGND VGND VPWR VPWR _13694_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12645_ _12645_/A _12645_/B VGND VGND VPWR VPWR _12645_/X sky130_fd_sc_hd__or2_1
XFILLER_157_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12576_ _12570_/Y _12619_/A _12614_/A _14740_/Q _12575_/X VGND VGND VPWR VPWR _12576_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_129_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14315_ _14617_/CLK _14315_/D VGND VGND VPWR VPWR _14315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11527_ _13624_/Q _11529_/B VGND VGND VPWR VPWR _11528_/A sky130_fd_sc_hd__and2_1
XFILLER_144_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold309 hold309/A VGND VGND VPWR VPWR hold309/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14246_ _14256_/CLK _14246_/D VGND VGND VPWR VPWR _14246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11458_ _11458_/A VGND VGND VPWR VPWR _13821_/D sky130_fd_sc_hd__clkbuf_1
X_10409_ _10396_/X _10400_/B _10397_/A VGND VGND VPWR VPWR _10410_/B sky130_fd_sc_hd__a21oi_1
XFILLER_124_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14177_ _14196_/CLK _14177_/D VGND VGND VPWR VPWR _14177_/Q sky130_fd_sc_hd__dfxtp_1
X_11389_ _11389_/A VGND VGND VPWR VPWR _13787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14760__71 VGND VGND VPWR VPWR _14760__71/HI _13387_/D sky130_fd_sc_hd__conb_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _14588_/CLK _14631_/Q VGND VGND VPWR VPWR hold212/A sky130_fd_sc_hd__dfxtp_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05950_ _05950_/A _05950_/B _05950_/C VGND VGND VPWR VPWR _05951_/D sky130_fd_sc_hd__and3_1
X_13059_ _13562_/CLK _13059_/D VGND VGND VPWR VPWR hold320/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07620_ _07620_/A _07620_/B VGND VGND VPWR VPWR _07635_/A sky130_fd_sc_hd__and2_1
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07551_ _07556_/A _07551_/B VGND VGND VPWR VPWR _07559_/A sky130_fd_sc_hd__nand2_1
XFILLER_35_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06502_ _06502_/A _10349_/A _06504_/B VGND VGND VPWR VPWR _06505_/B sky130_fd_sc_hd__and3_1
XFILLER_62_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07482_ _13148_/Q _09206_/B VGND VGND VPWR VPWR _07483_/B sky130_fd_sc_hd__or2_1
XFILLER_50_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09221_ _13539_/Q _13540_/Q _13541_/Q _13542_/Q _09250_/B VGND VGND VPWR VPWR _09244_/A
+ sky130_fd_sc_hd__o41a_1
X_06433_ _06433_/A _06433_/B VGND VGND VPWR VPWR _06437_/A sky130_fd_sc_hd__nand2_1
XFILLER_148_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09152_ _09153_/B _09153_/C _13534_/Q VGND VGND VPWR VPWR _09159_/B sky130_fd_sc_hd__a21oi_1
X_06364_ _06363_/Y _06030_/B _14633_/D _14640_/Q VGND VGND VPWR VPWR _14429_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_148_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08103_ _13426_/Q VGND VGND VPWR VPWR _08162_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06295_ _14162_/Q _14206_/D VGND VGND VPWR VPWR _06295_/Y sky130_fd_sc_hd__nor2_1
X_09083_ _09083_/A VGND VGND VPWR VPWR _12774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08034_ _12955_/Q _13255_/Q _08040_/S VGND VGND VPWR VPWR _08035_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09985_ _09984_/X _09977_/X _10596_/B VGND VGND VPWR VPWR _09986_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08936_ _08903_/A _08903_/B _08909_/A _08909_/B VGND VGND VPWR VPWR _08963_/B sky130_fd_sc_hd__a22o_1
XFILLER_57_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08867_ _08944_/A _08867_/B VGND VGND VPWR VPWR _08867_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_111_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07818_ _13255_/Q _07819_/B VGND VGND VPWR VPWR _07833_/A sky130_fd_sc_hd__nor2_1
XFILLER_57_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08798_ _08851_/A VGND VGND VPWR VPWR _08828_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07749_ _07724_/A _07726_/B _07724_/B VGND VGND VPWR VPWR _07750_/A sky130_fd_sc_hd__o21ba_1
XFILLER_25_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10760_ _13002_/Q _10768_/B VGND VGND VPWR VPWR _10761_/A sky130_fd_sc_hd__and2_1
XFILLER_53_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09419_ _09419_/A _09419_/B _09419_/C _09419_/D VGND VGND VPWR VPWR _09420_/D sky130_fd_sc_hd__nor4_2
XFILLER_158_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10691_ _10691_/A VGND VGND VPWR VPWR _12924_/D sky130_fd_sc_hd__clkbuf_1
X_12430_ _12480_/S VGND VGND VPWR VPWR _12439_/S sky130_fd_sc_hd__buf_2
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12361_ _12361_/A VGND VGND VPWR VPWR _14603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14100_ _14319_/CLK _14100_/D VGND VGND VPWR VPWR _14100_/Q sky130_fd_sc_hd__dfxtp_1
X_11312_ _11312_/A VGND VGND VPWR VPWR _13764_/D sky130_fd_sc_hd__clkbuf_1
X_12292_ _12292_/A VGND VGND VPWR VPWR _14562_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14031_ _14721_/CLK _14031_/D VGND VGND VPWR VPWR _14031_/Q sky130_fd_sc_hd__dfxtp_1
X_11243_ _13339_/Q _10962_/A _11236_/X _11242_/Y VGND VGND VPWR VPWR _13339_/D sky130_fd_sc_hd__o22a_1
XFILLER_153_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11174_ _14612_/Q _14574_/Q _14505_/Q _14457_/Q _11115_/X _11116_/X VGND VGND VPWR
+ VPWR _11175_/A sky130_fd_sc_hd__mux4_1
XFILLER_161_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10125_ _13863_/Q _13847_/Q _14167_/D VGND VGND VPWR VPWR _10126_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10056_ _10056_/A VGND VGND VPWR VPWR _10056_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13815_ _14633_/CLK hold324/X VGND VGND VPWR VPWR _13815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13746_ _14588_/CLK _13746_/D VGND VGND VPWR VPWR _13746_/Q sky130_fd_sc_hd__dfxtp_4
X_10958_ _12590_/A VGND VGND VPWR VPWR _10960_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13677_ _13681_/CLK _13677_/D repeater56/X VGND VGND VPWR VPWR _13677_/Q sky130_fd_sc_hd__dfrtp_1
X_10889_ _13161_/Q _10891_/B VGND VGND VPWR VPWR _10890_/A sky130_fd_sc_hd__and2_1
XFILLER_148_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12628_ _14741_/Q VGND VGND VPWR VPWR _12631_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12559_ _12559_/A VGND VGND VPWR VPWR _14724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06080_ _06256_/S VGND VGND VPWR VPWR _10023_/A sky130_fd_sc_hd__clkbuf_2
Xhold106 hold106/A VGND VGND VPWR VPWR hold106/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold117 hold117/A VGND VGND VPWR VPWR hold117/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold128 hold128/A VGND VGND VPWR VPWR hold128/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_99_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14229_ _14539_/CLK _14229_/D VGND VGND VPWR VPWR _14229_/Q sky130_fd_sc_hd__dfxtp_1
Xhold139 hold139/A VGND VGND VPWR VPWR hold139/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _09770_/A _09770_/B VGND VGND VPWR VPWR _09781_/A sky130_fd_sc_hd__or2_1
XFILLER_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06982_ _13022_/Q _13023_/Q _13024_/Q _13025_/Q _08002_/B VGND VGND VPWR VPWR _06982_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _13456_/Q _08746_/A VGND VGND VPWR VPWR _08724_/A sky130_fd_sc_hd__nand2_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05933_ _13720_/Q _13729_/Q _13730_/Q _13731_/Q VGND VGND VPWR VPWR _05934_/C sky130_fd_sc_hd__or4_1
XFILLER_66_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08652_ _08653_/A _08654_/A _08653_/B VGND VGND VPWR VPWR _08652_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_54_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07603_ _13746_/Q _13106_/Q VGND VGND VPWR VPWR _07800_/S sky130_fd_sc_hd__xor2_4
XFILLER_26_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08583_ _08607_/A VGND VGND VPWR VPWR _08591_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07534_ _13151_/Q _13152_/Q _13153_/Q _13154_/Q _09257_/B VGND VGND VPWR VPWR _07534_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07465_ _07477_/B _07504_/A VGND VGND VPWR VPWR _07465_/Y sky130_fd_sc_hd__xnor2_1
X_09204_ _09182_/X _09202_/X _09203_/Y _07575_/X VGND VGND VPWR VPWR _13540_/D sky130_fd_sc_hd__a31o_1
X_06416_ _06469_/A hold187/A _06455_/A VGND VGND VPWR VPWR _06416_/X sky130_fd_sc_hd__and3b_1
XFILLER_50_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07396_ _07396_/A _09151_/B VGND VGND VPWR VPWR _07396_/X sky130_fd_sc_hd__and2_1
X_09135_ _09135_/A _09135_/B _09135_/C VGND VGND VPWR VPWR _09137_/B sky130_fd_sc_hd__and3_1
X_06347_ hold77/A _14401_/D _14402_/D _14405_/D VGND VGND VPWR VPWR _06348_/D sky130_fd_sc_hd__and4_1
XFILLER_163_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09066_ _09600_/A VGND VGND VPWR VPWR _09075_/S sky130_fd_sc_hd__clkbuf_2
X_06278_ _06278_/A VGND VGND VPWR VPWR _13957_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08017_ _08018_/B _08018_/C _08018_/A VGND VGND VPWR VPWR _08017_/X sky130_fd_sc_hd__a21o_1
XFILLER_118_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09968_ _13507_/Q _13696_/Q _09968_/S VGND VGND VPWR VPWR _09969_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08919_ _08919_/A _08919_/B VGND VGND VPWR VPWR _08919_/Y sky130_fd_sc_hd__nor2_1
XFILLER_58_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09899_ _13697_/Q _13698_/Q _09886_/A _09893_/B _09672_/Y VGND VGND VPWR VPWR _09899_/X
+ sky130_fd_sc_hd__a41o_1
X_11930_ _11930_/A VGND VGND VPWR VPWR _14271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _11861_/A VGND VGND VPWR VPWR _14228_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _13621_/CLK _13600_/D repeater56/X VGND VGND VPWR VPWR _13600_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10812_ _13026_/Q _10812_/B VGND VGND VPWR VPWR _10813_/A sky130_fd_sc_hd__and2_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _14619_/CLK _14580_/D VGND VGND VPWR VPWR _14580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11792_ _11792_/A VGND VGND VPWR VPWR _14089_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13531_ _13532_/CLK _13531_/D hold1/X VGND VGND VPWR VPWR _13531_/Q sky130_fd_sc_hd__dfrtp_2
X_10743_ _10743_/A VGND VGND VPWR VPWR _12948_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13462_ _13855_/CLK _13462_/D repeater57/X VGND VGND VPWR VPWR _13462_/Q sky130_fd_sc_hd__dfrtp_1
X_10674_ _10674_/A VGND VGND VPWR VPWR _12917_/D sky130_fd_sc_hd__clkbuf_1
X_12413_ _12413_/A VGND VGND VPWR VPWR _14640_/D sky130_fd_sc_hd__clkbuf_1
X_13393_ _13593_/CLK hold399/X VGND VGND VPWR VPWR _13393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12344_ _12394_/S VGND VGND VPWR VPWR _12353_/S sky130_fd_sc_hd__buf_2
XFILLER_5_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12275_ _12275_/A VGND VGND VPWR VPWR _14552_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14014_ _14533_/CLK _14014_/D VGND VGND VPWR VPWR _14014_/Q sky130_fd_sc_hd__dfxtp_1
X_11226_ _14616_/Q _14578_/Q _14509_/Q _14461_/Q _11186_/X _11187_/X VGND VGND VPWR
+ VPWR _11227_/A sky130_fd_sc_hd__mux4_1
XFILLER_122_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11157_ _11224_/A VGND VGND VPWR VPWR _11157_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10108_ _14143_/D _14210_/Q _14142_/D _06117_/X _14208_/Q VGND VGND VPWR VPWR _14156_/D
+ sky130_fd_sc_hd__a221o_1
X_11088_ _11207_/A VGND VGND VPWR VPWR _11088_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10039_ _10039_/A VGND VGND VPWR VPWR _13945_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13729_ _13805_/CLK hold303/X VGND VGND VPWR VPWR _13729_/Q sky130_fd_sc_hd__dfxtp_1
X_07250_ _09086_/B VGND VGND VPWR VPWR _07261_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06201_ _06200_/X _06196_/X _10193_/A VGND VGND VPWR VPWR _06202_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07181_ _07182_/A _07182_/B _07182_/C VGND VGND VPWR VPWR _07183_/A sky130_fd_sc_hd__a21oi_1
XFILLER_8_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06132_ _06132_/A VGND VGND VPWR VPWR _14151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06063_ _13973_/Q _13971_/Q _10020_/A VGND VGND VPWR VPWR _06063_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09822_ _09822_/A _09822_/B VGND VGND VPWR VPWR _09824_/A sky130_fd_sc_hd__nor2_1
XFILLER_101_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09753_ _09753_/A _09753_/B VGND VGND VPWR VPWR _09753_/X sky130_fd_sc_hd__xor2_1
XFILLER_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06965_ _06874_/X _06964_/X _06897_/X VGND VGND VPWR VPWR _13023_/D sky130_fd_sc_hd__a21o_1
XFILLER_67_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08704_ _08704_/A _08704_/B _08714_/C VGND VGND VPWR VPWR _08704_/Y sky130_fd_sc_hd__nand3_1
XFILLER_104_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05916_ _13726_/Q _13727_/Q _13728_/Q _13733_/Q VGND VGND VPWR VPWR _05917_/D sky130_fd_sc_hd__and4_1
XFILLER_27_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09684_ _09778_/B _09672_/Y _09679_/C _09683_/X VGND VGND VPWR VPWR _13668_/D sky130_fd_sc_hd__a31o_1
XFILLER_66_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06896_ _07940_/A VGND VGND VPWR VPWR _07932_/A sky130_fd_sc_hd__buf_2
XFILLER_27_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08635_ _08645_/A _08635_/B VGND VGND VPWR VPWR _08635_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ _08581_/A _08566_/B VGND VGND VPWR VPWR _08567_/C sky130_fd_sc_hd__and2_1
XFILLER_120_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07517_ _07519_/A _07532_/B VGND VGND VPWR VPWR _07517_/Y sky130_fd_sc_hd__nand2_1
X_08497_ _08521_/A _08497_/B _13438_/Q VGND VGND VPWR VPWR _08497_/Y sky130_fd_sc_hd__nand3b_1
X_07448_ _07400_/A _07345_/X _07420_/A VGND VGND VPWR VPWR _07450_/A sky130_fd_sc_hd__o21a_1
XFILLER_22_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07379_ _13140_/Q _09139_/B _09139_/C VGND VGND VPWR VPWR _07381_/A sky130_fd_sc_hd__and3_1
XFILLER_129_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09118_ _13529_/Q _09118_/B VGND VGND VPWR VPWR _09134_/C sky130_fd_sc_hd__xnor2_1
XFILLER_164_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10390_ _10390_/A _10390_/B VGND VGND VPWR VPWR _10391_/B sky130_fd_sc_hd__nor2_1
XFILLER_89_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09049_ _13224_/Q _13453_/Q _09051_/S VGND VGND VPWR VPWR _09050_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12060_ _12060_/A VGND VGND VPWR VPWR _14448_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold470 hold470/A VGND VGND VPWR VPWR hold470/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold481 hold481/A VGND VGND VPWR VPWR hold481/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_11011_ _11163_/A VGND VGND VPWR VPWR _11011_/X sky130_fd_sc_hd__buf_2
Xhold492 hold492/A VGND VGND VPWR VPWR hold492/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12962_ _13263_/CLK hold107/X VGND VGND VPWR VPWR _12962_/Q sky130_fd_sc_hd__dfxtp_1
X_11913_ _11913_/A VGND VGND VPWR VPWR _14263_/D sky130_fd_sc_hd__clkbuf_1
X_14701_ _14710_/CLK hold309/X VGND VGND VPWR VPWR _14701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12893_ _12970_/CLK _12893_/D hold1/X VGND VGND VPWR VPWR _12893_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _14644_/CLK _14645_/Q VGND VGND VPWR VPWR _14632_/Q sky130_fd_sc_hd__dfxtp_1
X_11844_ _11894_/S VGND VGND VPWR VPWR _11853_/S sky130_fd_sc_hd__buf_2
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _14712_/CLK _14563_/D VGND VGND VPWR VPWR _14563_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _11834_/B VGND VGND VPWR VPWR _11784_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_158_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10726_ _10726_/A VGND VGND VPWR VPWR _12940_/D sky130_fd_sc_hd__clkbuf_1
X_13514_ _14010_/CLK _13514_/D VGND VGND VPWR VPWR _13703_/D sky130_fd_sc_hd__dfxtp_1
X_14494_ _14495_/CLK _14494_/D VGND VGND VPWR VPWR _14494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13445_ _13598_/CLK _13445_/D repeater56/X VGND VGND VPWR VPWR _13445_/Q sky130_fd_sc_hd__dfrtp_1
X_10657_ _14337_/Q _14334_/Q _10656_/X VGND VGND VPWR VPWR _10657_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_139_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13376_ _14530_/CLK _13376_/D _12609_/A VGND VGND VPWR VPWR _13376_/Q sky130_fd_sc_hd__dfrtp_1
X_10588_ _10588_/A VGND VGND VPWR VPWR _13472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12327_ _12327_/A VGND VGND VPWR VPWR _14578_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12258_ _12258_/A VGND VGND VPWR VPWR _14544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11209_ _11209_/A VGND VGND VPWR VPWR _11209_/X sky130_fd_sc_hd__buf_2
XFILLER_122_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12189_ _12189_/A VGND VGND VPWR VPWR _14505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06750_ _13351_/Q _13347_/Q _13349_/Q _13345_/Q _13038_/Q _06746_/S VGND VGND VPWR
+ VPWR _06751_/B sky130_fd_sc_hd__mux4_1
X_06681_ _06681_/A _06681_/B _06681_/C VGND VGND VPWR VPWR _06681_/X sky130_fd_sc_hd__or3_1
XFILLER_37_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08420_ _09323_/A VGND VGND VPWR VPWR _09299_/S sky130_fd_sc_hd__buf_2
XFILLER_24_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08351_ _08351_/A VGND VGND VPWR VPWR _12710_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07302_ _09099_/A _07302_/B VGND VGND VPWR VPWR _09113_/B sky130_fd_sc_hd__xor2_4
XFILLER_32_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08282_ _08282_/A _08282_/B VGND VGND VPWR VPWR _08285_/A sky130_fd_sc_hd__nor2_1
X_07233_ _07461_/B _07249_/C VGND VGND VPWR VPWR _09088_/B sky130_fd_sc_hd__xor2_4
XFILLER_137_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07164_ _07164_/A _07164_/B VGND VGND VPWR VPWR _07166_/A sky130_fd_sc_hd__nor2_1
XFILLER_157_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06115_ _06115_/A VGND VGND VPWR VPWR _13963_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07095_ _07107_/A _07095_/B VGND VGND VPWR VPWR _07126_/B sky130_fd_sc_hd__xnor2_1
XFILLER_161_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06046_ _13969_/Q _13967_/Q _13977_/Q VGND VGND VPWR VPWR _06046_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09805_ _09795_/A _09804_/Y _09795_/B _09792_/A VGND VGND VPWR VPWR _09806_/B sky130_fd_sc_hd__a31o_1
XFILLER_59_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07997_ _06976_/X _07996_/Y _07932_/X VGND VGND VPWR VPWR _13279_/D sky130_fd_sc_hd__a21o_1
XFILLER_75_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06948_ _06948_/A _06948_/B _06950_/B VGND VGND VPWR VPWR _06948_/X sky130_fd_sc_hd__or3_1
X_09736_ _09736_/A VGND VGND VPWR VPWR _09778_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09667_ _09767_/A _09768_/B _09664_/X _09704_/A VGND VGND VPWR VPWR _09678_/C sky130_fd_sc_hd__a22o_1
XFILLER_43_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06879_ _06846_/A _06877_/A _06876_/A _06876_/B VGND VGND VPWR VPWR _06879_/X sky130_fd_sc_hd__a211o_1
XFILLER_28_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ _13445_/Q _09438_/B _08620_/B VGND VGND VPWR VPWR _08618_/X sky130_fd_sc_hd__a21o_1
XFILLER_27_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _13397_/Q _13595_/Q _09598_/S VGND VGND VPWR VPWR _09599_/A sky130_fd_sc_hd__mux2_2
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _14254_/Q _14250_/Q _14252_/Q _14248_/Q _13475_/Q _08545_/S VGND VGND VPWR
+ VPWR _08550_/B sky130_fd_sc_hd__mux4_1
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11560_ _11560_/A VGND VGND VPWR VPWR _13862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10511_ _10521_/B _14431_/D VGND VGND VPWR VPWR _10511_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11491_ _14518_/Q VGND VGND VPWR VPWR _11491_/X sky130_fd_sc_hd__buf_2
XFILLER_149_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13230_ _13617_/CLK hold411/X VGND VGND VPWR VPWR _13230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10442_ _10439_/Y _10439_/A _10449_/A VGND VGND VPWR VPWR _10443_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13161_ _13554_/CLK _13161_/D _12609_/A VGND VGND VPWR VPWR _13161_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10373_ _13519_/Q VGND VGND VPWR VPWR _10423_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_3_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12112_ _12112_/A VGND VGND VPWR VPWR _14471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13092_ _13562_/CLK hold320/X VGND VGND VPWR VPWR _13092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12043_ _12093_/S VGND VGND VPWR VPWR _12052_/S sky130_fd_sc_hd__buf_2
XFILLER_78_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13994_ _14720_/CLK _13994_/D VGND VGND VPWR VPWR _13994_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12945_ _13280_/CLK _12945_/D VGND VGND VPWR VPWR hold256/A sky130_fd_sc_hd__dfxtp_1
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _12881_/CLK _12876_/D hold1/X VGND VGND VPWR VPWR _12876_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14615_ _14615_/CLK _14615_/D VGND VGND VPWR VPWR _14615_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _11827_/A VGND VGND VPWR VPWR _14105_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _11354_/X _14070_/Q _11758_/S VGND VGND VPWR VPWR _11759_/A sky130_fd_sc_hd__mux2_1
X_14546_ _14720_/CLK _14546_/D VGND VGND VPWR VPWR _14546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10709_ _12890_/Q _10709_/B VGND VGND VPWR VPWR _10710_/A sky130_fd_sc_hd__and2_1
X_14477_ _14602_/CLK _14477_/D VGND VGND VPWR VPWR _14477_/Q sky130_fd_sc_hd__dfxtp_1
X_11689_ _14027_/Q _11494_/X _11689_/S VGND VGND VPWR VPWR _11690_/A sky130_fd_sc_hd__mux2_1
X_13428_ _14687_/CLK hold186/X VGND VGND VPWR VPWR _13428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13359_ _13359_/CLK _13359_/D hold1/X VGND VGND VPWR VPWR _13359_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07920_ _07914_/A _07912_/B _07917_/Y _07898_/B _07919_/Y VGND VGND VPWR VPWR _07925_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_111_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07851_ _06757_/B _07850_/Y _07861_/S VGND VGND VPWR VPWR _07852_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06802_ _13008_/Q _06807_/A VGND VGND VPWR VPWR _06825_/A sky130_fd_sc_hd__xnor2_1
X_07782_ _07782_/A VGND VGND VPWR VPWR _13663_/D sky130_fd_sc_hd__clkbuf_1
Xinput2 data_i[10] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09521_ _09513_/A _09514_/X _09534_/B _08733_/X VGND VGND VPWR VPWR _09521_/X sky130_fd_sc_hd__a31o_1
XFILLER_83_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06733_ _06871_/A _06733_/B _06737_/A VGND VGND VPWR VPWR _06733_/X sky130_fd_sc_hd__and3_1
XFILLER_65_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09452_ _09460_/A _09452_/B VGND VGND VPWR VPWR _09455_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06664_ _06664_/A VGND VGND VPWR VPWR _12999_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08403_ _08403_/A VGND VGND VPWR VPWR _12733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09383_ _13591_/Q _09383_/B VGND VGND VPWR VPWR _09383_/X sky130_fd_sc_hd__and2_1
X_06595_ _12898_/Q _06595_/B _06598_/D VGND VGND VPWR VPWR _06597_/A sky130_fd_sc_hd__and3_1
X_08334_ _13382_/Q _08333_/A _08298_/X VGND VGND VPWR VPWR _08334_/Y sky130_fd_sc_hd__o21ai_1
X_08265_ _08265_/A _08265_/B VGND VGND VPWR VPWR _08267_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07216_ _07209_/Y _07215_/Y _07218_/S VGND VGND VPWR VPWR _07217_/A sky130_fd_sc_hd__mux2_1
X_08196_ _08114_/X _08141_/X _08147_/B _08162_/Y VGND VGND VPWR VPWR _08199_/B sky130_fd_sc_hd__o22a_1
XFILLER_146_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07147_ _07147_/A _07147_/B VGND VGND VPWR VPWR _07149_/A sky130_fd_sc_hd__xor2_2
XFILLER_133_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07078_ _07101_/A _07078_/B VGND VGND VPWR VPWR _07079_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06029_ _14645_/Q _14641_/Q _14642_/Q _14643_/Q VGND VGND VPWR VPWR _06030_/B sky130_fd_sc_hd__and4_1
XFILLER_0_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09719_ _09717_/X _09673_/X _09718_/Y _09664_/X VGND VGND VPWR VPWR _09720_/C sky130_fd_sc_hd__o22a_1
X_10991_ _11262_/A VGND VGND VPWR VPWR _10991_/X sky130_fd_sc_hd__buf_2
XFILLER_16_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _13617_/CLK _12730_/D VGND VGND VPWR VPWR hold443/A sky130_fd_sc_hd__dfxtp_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _14737_/CLK _12661_/D _12609_/A VGND VGND VPWR VPWR _12662_/D sky130_fd_sc_hd__dfrtp_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11612_ _13983_/Q _11462_/X _11612_/S VGND VGND VPWR VPWR _11613_/A sky130_fd_sc_hd__mux2_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _14410_/CLK _14400_/D VGND VGND VPWR VPWR _14400_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _10901_/A _10900_/Y _11185_/A _12591_/X VGND VGND VPWR VPWR _12592_/X sky130_fd_sc_hd__o22a_1
X_11543_ _11591_/B VGND VGND VPWR VPWR _11552_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14331_ _14696_/CLK hold78/X VGND VGND VPWR VPWR hold432/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14262_ _14710_/CLK _14262_/D VGND VGND VPWR VPWR _14262_/Q sky130_fd_sc_hd__dfxtp_1
X_11474_ _11474_/A VGND VGND VPWR VPWR _13826_/D sky130_fd_sc_hd__clkbuf_1
X_13213_ _13598_/CLK _13213_/D VGND VGND VPWR VPWR _13213_/Q sky130_fd_sc_hd__dfxtp_1
X_10425_ _10426_/A _10426_/B _10426_/C VGND VGND VPWR VPWR _10431_/B sky130_fd_sc_hd__o21ai_1
X_14193_ _14693_/CLK _14193_/D VGND VGND VPWR VPWR _14194_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_124_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13144_ _13535_/CLK _13144_/D repeater57/X VGND VGND VPWR VPWR _13144_/Q sky130_fd_sc_hd__dfrtp_1
X_10356_ _13780_/Q _13781_/Q VGND VGND VPWR VPWR _10357_/B sky130_fd_sc_hd__and2_1
XFILLER_151_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13075_ _13076_/CLK _13075_/D VGND VGND VPWR VPWR _13075_/Q sky130_fd_sc_hd__dfxtp_1
X_10287_ _10287_/A VGND VGND VPWR VPWR _12666_/D sky130_fd_sc_hd__clkbuf_1
X_12026_ _14318_/Q _12025_/X _12026_/S VGND VGND VPWR VPWR _12027_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13977_ _14179_/CLK _13977_/D VGND VGND VPWR VPWR _13977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12928_ _13263_/CLK _12928_/D VGND VGND VPWR VPWR hold261/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _13805_/CLK _12859_/D VGND VGND VPWR VPWR hold319/A sky130_fd_sc_hd__dfxtp_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06380_ _14439_/Q _14437_/Q _14435_/Q _14433_/Q _13106_/D _13107_/D VGND VGND VPWR
+ VPWR _06495_/C sky130_fd_sc_hd__mux4_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14529_ _14555_/CLK _14529_/D VGND VGND VPWR VPWR hold132/A sky130_fd_sc_hd__dfxtp_1
XFILLER_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08050_ _08050_/A VGND VGND VPWR VPWR _12686_/D sky130_fd_sc_hd__clkbuf_1
X_07001_ _07001_/A _07001_/B _07001_/C VGND VGND VPWR VPWR _07001_/Y sky130_fd_sc_hd__nand3_1
XFILLER_127_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08952_ _08952_/A _08952_/B VGND VGND VPWR VPWR _08954_/A sky130_fd_sc_hd__nor2_1
XFILLER_69_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07903_ _07914_/A _07903_/B VGND VGND VPWR VPWR _07916_/A sky130_fd_sc_hd__nand2_1
X_08883_ _08895_/A _08883_/B VGND VGND VPWR VPWR _08914_/B sky130_fd_sc_hd__xnor2_1
XFILLER_97_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07834_ _13257_/Q _07840_/B VGND VGND VPWR VPWR _07858_/B sky130_fd_sc_hd__xnor2_2
XFILLER_56_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07765_ _07765_/A _07765_/B VGND VGND VPWR VPWR _07766_/B sky130_fd_sc_hd__nor2_1
XFILLER_44_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09504_ _09505_/A _09505_/B _09509_/D VGND VGND VPWR VPWR _09504_/X sky130_fd_sc_hd__a21o_1
X_06716_ _06716_/A VGND VGND VPWR VPWR _06716_/Y sky130_fd_sc_hd__inv_2
X_07696_ _07696_/A _07696_/B VGND VGND VPWR VPWR _07697_/B sky130_fd_sc_hd__or2_1
XFILLER_52_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09435_ _09454_/A _09454_/C _09454_/B VGND VGND VPWR VPWR _09435_/Y sky130_fd_sc_hd__o21ai_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06647_ _13037_/Q VGND VGND VPWR VPWR _06705_/S sky130_fd_sc_hd__clkbuf_2
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09366_ _09370_/B _09366_/B VGND VGND VPWR VPWR _13589_/D sky130_fd_sc_hd__xnor2_1
X_06578_ _12892_/Q _06574_/X _12893_/Q VGND VGND VPWR VPWR _06578_/Y sky130_fd_sc_hd__a21oi_1
X_08317_ _13376_/Q _13377_/Q _08317_/C _08317_/D VGND VGND VPWR VPWR _08325_/D sky130_fd_sc_hd__and4_1
XFILLER_138_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_40 _13333_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09297_ _13287_/Q _13525_/Q _09299_/S VGND VGND VPWR VPWR _09298_/A sky130_fd_sc_hd__mux2_1
XANTENNA_51 hold499/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 hold159/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_73 _10831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08248_ _08243_/B _08247_/Y _08286_/S VGND VGND VPWR VPWR _08249_/A sky130_fd_sc_hd__mux2_1
XANTENNA_84 input19/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_95 input12/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08179_ _08114_/X _08173_/X _08175_/X _08178_/Y VGND VGND VPWR VPWR _08180_/B sky130_fd_sc_hd__o211a_2
XFILLER_137_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10210_ _06215_/C _06216_/Y _10206_/S _10198_/X VGND VGND VPWR VPWR _14421_/D sky130_fd_sc_hd__o22a_1
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11190_ _11190_/A VGND VGND VPWR VPWR _11240_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10141_ _14282_/D _10149_/B VGND VGND VPWR VPWR _10147_/A sky130_fd_sc_hd__and2_1
XFILLER_0_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10072_ _14050_/D _13908_/D VGND VGND VPWR VPWR _10072_/X sky130_fd_sc_hd__and2_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13900_ _14209_/CLK hold441/X VGND VGND VPWR VPWR hold295/A sky130_fd_sc_hd__dfxtp_1
X_13831_ _14713_/CLK _13831_/D VGND VGND VPWR VPWR _13831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10974_ _11190_/A VGND VGND VPWR VPWR _11035_/A sky130_fd_sc_hd__buf_2
XFILLER_16_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13762_ _14710_/CLK _13762_/D VGND VGND VPWR VPWR _13762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12713_ _13596_/CLK _12713_/D VGND VGND VPWR VPWR hold377/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13693_ _13811_/CLK _13693_/D repeater57/X VGND VGND VPWR VPWR _13693_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_70_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12644_ _12631_/B _12567_/X _12643_/X _12617_/X VGND VGND VPWR VPWR _14746_/D sky130_fd_sc_hd__o211a_1
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12575_ _12573_/Y _11655_/A _14739_/Q _12568_/Y VGND VGND VPWR VPWR _12575_/X sky130_fd_sc_hd__a2bb2o_1
X_14314_ _14510_/CLK _14314_/D VGND VGND VPWR VPWR _14314_/Q sky130_fd_sc_hd__dfxtp_1
X_11526_ _11526_/A VGND VGND VPWR VPWR _13847_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11457_ _13821_/Q _11456_/X _11463_/S VGND VGND VPWR VPWR _11458_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14245_ _14256_/CLK _14245_/D VGND VGND VPWR VPWR _14245_/Q sky130_fd_sc_hd__dfxtp_1
X_10408_ _10421_/A _10411_/C VGND VGND VPWR VPWR _10410_/A sky130_fd_sc_hd__and2b_1
X_14176_ _14196_/CLK _14176_/D VGND VGND VPWR VPWR _14176_/Q sky130_fd_sc_hd__dfxtp_1
X_11388_ _13718_/Q _11394_/B VGND VGND VPWR VPWR _11389_/A sky130_fd_sc_hd__and2_1
XFILLER_125_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13127_ _14645_/CLK _14630_/Q VGND VGND VPWR VPWR hold62/A sky130_fd_sc_hd__dfxtp_2
XFILLER_113_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10339_ _10339_/A hold131/A _10339_/C VGND VGND VPWR VPWR _10340_/B sky130_fd_sc_hd__nor3_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _13562_/CLK _13058_/D VGND VGND VPWR VPWR hold310/A sky130_fd_sc_hd__dfxtp_1
XFILLER_140_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12009_ _12009_/A VGND VGND VPWR VPWR _14312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07550_ _13157_/Q _09258_/B VGND VGND VPWR VPWR _07551_/B sky130_fd_sc_hd__or2_1
XFILLER_19_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06501_ _06500_/A _06498_/X _06499_/Y _06500_/Y VGND VGND VPWR VPWR _12884_/D sky130_fd_sc_hd__o31ai_1
XFILLER_34_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07481_ _07481_/A VGND VGND VPWR VPWR _09206_/B sky130_fd_sc_hd__clkbuf_2
X_09220_ _09220_/A _09220_/B _09220_/C _09220_/D VGND VGND VPWR VPWR _09242_/B sky130_fd_sc_hd__or4_1
XFILLER_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06432_ _12879_/Q _06450_/B VGND VGND VPWR VPWR _06433_/B sky130_fd_sc_hd__nand2_1
X_09151_ _13533_/Q _09151_/B VGND VGND VPWR VPWR _09156_/A sky130_fd_sc_hd__nand2_1
X_06363_ _14644_/Q VGND VGND VPWR VPWR _06363_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_147_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08102_ _08199_/A VGND VGND VPWR VPWR _08220_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_09082_ _13238_/Q _13467_/Q _09587_/S VGND VGND VPWR VPWR _09083_/A sky130_fd_sc_hd__mux2_1
X_06294_ _06292_/A _06292_/Y _14197_/D _06293_/X VGND VGND VPWR VPWR _14207_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08033_ _08033_/A VGND VGND VPWR VPWR _12675_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09984_ _14593_/Q _14591_/Q _10597_/A VGND VGND VPWR VPWR _09984_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08935_ _08935_/A _08935_/B VGND VGND VPWR VPWR _08937_/A sky130_fd_sc_hd__xor2_1
XFILLER_130_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08866_ _08889_/A _08866_/B VGND VGND VPWR VPWR _08867_/B sky130_fd_sc_hd__nand2_1
XFILLER_96_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07817_ _07811_/X _07815_/Y _07816_/X _06685_/X VGND VGND VPWR VPWR _13254_/D sky130_fd_sc_hd__a31o_1
X_08797_ _14003_/Q VGND VGND VPWR VPWR _08851_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07748_ _07748_/A _07748_/B VGND VGND VPWR VPWR _07787_/A sky130_fd_sc_hd__xnor2_1
XFILLER_37_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07679_ _07649_/A _07651_/B _07649_/B VGND VGND VPWR VPWR _07680_/B sky130_fd_sc_hd__o21ba_1
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09418_ _09396_/A _09400_/Y _09401_/Y _09419_/C _09419_/D VGND VGND VPWR VPWR _09420_/C
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_52_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10690_ _12881_/Q _10698_/B VGND VGND VPWR VPWR _10691_/A sky130_fd_sc_hd__and2_1
XFILLER_9_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09349_ _09349_/A VGND VGND VPWR VPWR _12800_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12360_ _14603_/Q _11975_/X _12364_/S VGND VGND VPWR VPWR _12361_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11311_ _13764_/Q _11310_/X _11311_/S VGND VGND VPWR VPWR _11312_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12291_ _14562_/Q _11965_/X _12291_/S VGND VGND VPWR VPWR _12292_/A sky130_fd_sc_hd__mux2_1
X_14030_ _14275_/CLK _14030_/D VGND VGND VPWR VPWR _14030_/Q sky130_fd_sc_hd__dfxtp_1
X_11242_ _11242_/A _11242_/B VGND VGND VPWR VPWR _11242_/Y sky130_fd_sc_hd__nand2_1
XFILLER_162_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11173_ _11136_/X _11170_/X _11172_/X _11157_/X VGND VGND VPWR VPWR _11173_/X sky130_fd_sc_hd__o211a_1
X_10124_ _06145_/D _06292_/Y _14197_/D _10116_/X VGND VGND VPWR VPWR _14205_/D sky130_fd_sc_hd__a22o_1
XFILLER_164_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10055_ hold160/A _10056_/A _10060_/A VGND VGND VPWR VPWR _14039_/D sky130_fd_sc_hd__a21o_1
XFILLER_76_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13814_ _14647_/CLK _13814_/D VGND VGND VPWR VPWR _13814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13745_ _14179_/CLK hold228/X VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__dfxtp_1
X_10957_ _10957_/A VGND VGND VPWR VPWR _10957_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13676_ _13721_/CLK _13676_/D repeater56/X VGND VGND VPWR VPWR _13676_/Q sky130_fd_sc_hd__dfrtp_1
X_10888_ _10888_/A VGND VGND VPWR VPWR _13202_/D sky130_fd_sc_hd__clkbuf_1
X_12627_ _12631_/C _12626_/Y _12580_/X VGND VGND VPWR VPWR _14740_/D sky130_fd_sc_hd__o21ai_1
XFILLER_157_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12558_ _11365_/X _14724_/Q _12562_/S VGND VGND VPWR VPWR _12559_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11509_ _11509_/A VGND VGND VPWR VPWR _13837_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12489_ _12489_/A VGND VGND VPWR VPWR _14674_/D sky130_fd_sc_hd__clkbuf_1
Xhold107 hold107/A VGND VGND VPWR VPWR hold107/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold118 input24/X VGND VGND VPWR VPWR hold118/X sky130_fd_sc_hd__buf_8
Xhold129 hold129/A VGND VGND VPWR VPWR hold129/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_14228_ _14495_/CLK _14228_/D VGND VGND VPWR VPWR _14228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14159_ _14159_/CLK _14160_/Q VGND VGND VPWR VPWR hold272/A sky130_fd_sc_hd__dfxtp_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _06981_/A _06981_/B VGND VGND VPWR VPWR _06981_/Y sky130_fd_sc_hd__nor2_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05932_ _13732_/Q _13737_/Q _13738_/Q _13739_/Q VGND VGND VPWR VPWR _05934_/B sky130_fd_sc_hd__or4_1
X_08720_ _08741_/A _08718_/B _08713_/A VGND VGND VPWR VPWR _08728_/A sky130_fd_sc_hd__o21a_1
XFILLER_140_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08651_ _08664_/A _08651_/B VGND VGND VPWR VPWR _08653_/B sky130_fd_sc_hd__nand2_1
XFILLER_27_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07602_ _13169_/D _07602_/B VGND VGND VPWR VPWR _07602_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_54_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08582_ _08582_/A _08582_/B _08582_/C VGND VGND VPWR VPWR _08607_/A sky130_fd_sc_hd__nand3_1
XFILLER_35_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07533_ _07533_/A _07533_/B VGND VGND VPWR VPWR _07533_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07464_ _13147_/Q _07513_/B VGND VGND VPWR VPWR _07504_/A sky130_fd_sc_hd__xnor2_1
XFILLER_22_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09203_ _09205_/A _09220_/B VGND VGND VPWR VPWR _09203_/Y sky130_fd_sc_hd__nand2_1
X_06415_ _14433_/Q _14431_/Q _06425_/S VGND VGND VPWR VPWR _06415_/X sky130_fd_sc_hd__mux2_1
X_07395_ _07395_/A VGND VGND VPWR VPWR _09151_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_148_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09134_ _09134_/A _09134_/B _09134_/C _09134_/D VGND VGND VPWR VPWR _09135_/C sky130_fd_sc_hd__or4_1
XFILLER_148_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06346_ _06346_/A VGND VGND VPWR VPWR _14408_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09065_ _09065_/A VGND VGND VPWR VPWR _12766_/D sky130_fd_sc_hd__clkbuf_1
X_06277_ _13811_/Q _13795_/Q _06281_/S VGND VGND VPWR VPWR _06278_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08016_ _08016_/A _08016_/B VGND VGND VPWR VPWR _08018_/A sky130_fd_sc_hd__nand2_1
XFILLER_123_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09967_ _09967_/A VGND VGND VPWR VPWR _12869_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08918_ _08941_/A _08918_/B VGND VGND VPWR VPWR _08922_/B sky130_fd_sc_hd__or2_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _09896_/Y _09894_/C _09897_/X VGND VGND VPWR VPWR _13697_/D sky130_fd_sc_hd__a21oi_1
XFILLER_58_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08849_ _08929_/C VGND VGND VPWR VPWR _08978_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _14228_/Q _11472_/X _11864_/S VGND VGND VPWR VPWR _11861_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _10811_/A VGND VGND VPWR VPWR _13067_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ _13567_/Q _11795_/B VGND VGND VPWR VPWR _11792_/A sky130_fd_sc_hd__and2_1
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13530_ _13534_/CLK _13530_/D _12609_/A VGND VGND VPWR VPWR _13530_/Q sky130_fd_sc_hd__dfrtp_2
X_10742_ _12905_/Q _10742_/B VGND VGND VPWR VPWR _10743_/A sky130_fd_sc_hd__and2_1
XFILLER_41_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10673_ _10671_/X _10673_/B _10673_/C VGND VGND VPWR VPWR _10674_/A sky130_fd_sc_hd__and3b_1
X_13461_ _13626_/CLK _13461_/D repeater57/X VGND VGND VPWR VPWR _13461_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12412_ _12418_/A _12418_/B input26/X VGND VGND VPWR VPWR _12413_/A sky130_fd_sc_hd__and3_1
X_13392_ _14012_/CLK hold431/X VGND VGND VPWR VPWR _13392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12343_ _12377_/A VGND VGND VPWR VPWR _12394_/S sky130_fd_sc_hd__buf_2
X_12274_ _11365_/X _14552_/Q _12278_/S VGND VGND VPWR VPWR _12275_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11225_ _11207_/X _11221_/X _11223_/X _12647_/A VGND VGND VPWR VPWR _11225_/X sky130_fd_sc_hd__o211a_1
X_14013_ _14533_/CLK _14013_/D VGND VGND VPWR VPWR _14013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11156_ _11156_/A _11155_/X VGND VGND VPWR VPWR _11156_/X sky130_fd_sc_hd__or2b_1
XFILLER_122_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10107_ _10107_/A VGND VGND VPWR VPWR _14143_/D sky130_fd_sc_hd__inv_2
XFILLER_49_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11087_ _11065_/X _11080_/X _11085_/X _11086_/X VGND VGND VPWR VPWR _11087_/X sky130_fd_sc_hd__o211a_1
XFILLER_48_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10038_ _13799_/Q _13783_/Q _13935_/D VGND VGND VPWR VPWR _10039_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11989_ _14306_/Q _11988_/X _11998_/S VGND VGND VPWR VPWR _11990_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13728_ _13805_/CLK hold68/X VGND VGND VPWR VPWR _13728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13659_ _13666_/CLK _13659_/D VGND VGND VPWR VPWR _13659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06200_ _14421_/Q _14419_/Q _10194_/A VGND VGND VPWR VPWR _06200_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07180_ _07196_/A _07180_/B VGND VGND VPWR VPWR _07182_/C sky130_fd_sc_hd__nand2_1
XFILLER_145_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06131_ _06130_/X _06126_/X _10106_/A VGND VGND VPWR VPWR _06132_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06062_ _06062_/A VGND VGND VPWR VPWR _13919_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09821_ _13680_/Q _09821_/B VGND VGND VPWR VPWR _09822_/B sky130_fd_sc_hd__nor2_1
XFILLER_59_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09752_ _09725_/A _09726_/A _09725_/B _09741_/A _09751_/Y VGND VGND VPWR VPWR _09753_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_140_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06964_ _06967_/B _06964_/B VGND VGND VPWR VPWR _06964_/X sky130_fd_sc_hd__xor2_1
XFILLER_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08703_ _08704_/A _08704_/B _08714_/C VGND VGND VPWR VPWR _08709_/B sky130_fd_sc_hd__a21o_1
XFILLER_95_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05915_ _13722_/Q _13723_/Q _13724_/Q _13725_/Q VGND VGND VPWR VPWR _05915_/X sky130_fd_sc_hd__and4_1
XFILLER_66_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06895_ _06895_/A _06895_/B VGND VGND VPWR VPWR _07940_/A sky130_fd_sc_hd__and2_1
X_09683_ _09883_/B _09683_/B VGND VGND VPWR VPWR _09683_/X sky130_fd_sc_hd__and2_1
XFILLER_54_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08634_ _08634_/A VGND VGND VPWR VPWR _09457_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08565_ _08544_/X _08427_/A _08442_/A VGND VGND VPWR VPWR _08566_/B sky130_fd_sc_hd__o21a_1
XFILLER_54_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07516_ _07519_/A _07532_/B VGND VGND VPWR VPWR _07516_/X sky130_fd_sc_hd__or2_1
X_08496_ _08582_/A VGND VGND VPWR VPWR _08521_/A sky130_fd_sc_hd__buf_2
XFILLER_120_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07447_ _13145_/Q _09183_/B VGND VGND VPWR VPWR _07454_/A sky130_fd_sc_hd__nand2_1
XFILLER_149_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_170_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _14732_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07378_ _09139_/B _09139_/C VGND VGND VPWR VPWR _09140_/B sky130_fd_sc_hd__and2_1
XFILLER_129_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06329_ _06327_/Y _06328_/X _14424_/D VGND VGND VPWR VPWR _06330_/A sky130_fd_sc_hd__mux2_1
X_09117_ _09117_/A VGND VGND VPWR VPWR _13528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09048_ _09048_/A VGND VGND VPWR VPWR _12759_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold460 hold460/A VGND VGND VPWR VPWR hold460/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold471 hold471/A VGND VGND VPWR VPWR hold471/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_11010_ _12585_/A VGND VGND VPWR VPWR _11010_/X sky130_fd_sc_hd__buf_2
Xhold482 hold9/X VGND VGND VPWR VPWR hold482/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_78_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold493 hold493/A VGND VGND VPWR VPWR hold493/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_78_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12961_ _13263_/CLK hold261/X VGND VGND VPWR VPWR _12961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14700_ _14710_/CLK hold384/X VGND VGND VPWR VPWR _14700_/Q sky130_fd_sc_hd__dfxtp_1
X_11912_ _14263_/Q _11469_/X _11918_/S VGND VGND VPWR VPWR _11913_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _12970_/CLK _12892_/D hold1/X VGND VGND VPWR VPWR _12892_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _14679_/CLK hold205/X VGND VGND VPWR VPWR _14631_/Q sky130_fd_sc_hd__dfxtp_2
X_11843_ _11877_/A VGND VGND VPWR VPWR _11894_/S sky130_fd_sc_hd__buf_2
XFILLER_45_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _14600_/CLK _14562_/D VGND VGND VPWR VPWR _14562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _11819_/A VGND VGND VPWR VPWR _11834_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _14010_/CLK _13513_/D VGND VGND VPWR VPWR _13711_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_14_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10725_ _12897_/Q _10731_/B VGND VGND VPWR VPWR _10726_/A sky130_fd_sc_hd__and2_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14493_ _14598_/CLK _14493_/D VGND VGND VPWR VPWR _14493_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_161_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _14696_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13444_ _13702_/CLK _13444_/D repeater56/X VGND VGND VPWR VPWR _13444_/Q sky130_fd_sc_hd__dfrtp_1
X_10656_ _10673_/B VGND VGND VPWR VPWR _10656_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13375_ _13377_/CLK _13375_/D repeater57/X VGND VGND VPWR VPWR _13375_/Q sky130_fd_sc_hd__dfrtp_1
X_10587_ _13434_/Q hold504/A VGND VGND VPWR VPWR _10588_/A sky130_fd_sc_hd__or2_1
XFILLER_155_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12326_ _14578_/Q _12016_/X _12332_/S VGND VGND VPWR VPWR _12327_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12257_ _11323_/X _14544_/Q _12259_/S VGND VGND VPWR VPWR _12258_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11208_ _11208_/A VGND VGND VPWR VPWR _11208_/X sky130_fd_sc_hd__clkbuf_4
X_12188_ _14505_/Q _12004_/X _12194_/S VGND VGND VPWR VPWR _12189_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11139_ _14309_/Q _14479_/Q _14235_/Q _14065_/Q _11137_/X _11138_/X VGND VGND VPWR
+ VPWR _11139_/X sky130_fd_sc_hd__mux4_1
XFILLER_1_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06680_ _13000_/Q _07821_/B VGND VGND VPWR VPWR _06681_/C sky130_fd_sc_hd__and2_1
XFILLER_91_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08350_ _13074_/Q _13355_/Q _10891_/B VGND VGND VPWR VPWR _08351_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07301_ _07461_/A _07311_/B VGND VGND VPWR VPWR _07302_/B sky130_fd_sc_hd__and2_1
X_08281_ _13369_/Q _08281_/B VGND VGND VPWR VPWR _08282_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_152_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _14602_/CLK sky130_fd_sc_hd__clkbuf_16
X_07232_ _07266_/A _07227_/X _07228_/X _07361_/B _07231_/Y VGND VGND VPWR VPWR _07249_/C
+ sky130_fd_sc_hd__a32o_2
XFILLER_146_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07163_ _07163_/A _07163_/B _07163_/C VGND VGND VPWR VPWR _07164_/B sky130_fd_sc_hd__and3_1
XFILLER_9_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06114_ _13944_/D _06114_/B _06114_/C VGND VGND VPWR VPWR _06115_/A sky130_fd_sc_hd__or3_1
X_07094_ _07107_/B _07107_/C VGND VGND VPWR VPWR _07095_/B sky130_fd_sc_hd__nor2_1
XFILLER_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06045_ _12400_/C VGND VGND VPWR VPWR _14638_/D sky130_fd_sc_hd__inv_2
XFILLER_160_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09804_ _09804_/A VGND VGND VPWR VPWR _09804_/Y sky130_fd_sc_hd__inv_2
X_07996_ _07998_/B _07996_/B VGND VGND VPWR VPWR _07996_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09735_ _09735_/A VGND VGND VPWR VPWR _09836_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_28_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06947_ _06948_/A _06948_/B _06950_/B VGND VGND VPWR VPWR _06947_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09666_ _09718_/A _13711_/Q VGND VGND VPWR VPWR _09704_/A sky130_fd_sc_hd__and2b_1
X_06878_ _06870_/A _06868_/A _06868_/B VGND VGND VPWR VPWR _06878_/X sky130_fd_sc_hd__a21bo_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08617_ _09365_/A VGND VGND VPWR VPWR _08617_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09597_ _09597_/A VGND VGND VPWR VPWR _12813_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _13476_/Q VGND VGND VPWR VPWR _08578_/A sky130_fd_sc_hd__inv_2
XFILLER_70_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_143_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _14693_/CLK sky130_fd_sc_hd__clkbuf_16
X_08479_ _13437_/Q _09383_/B VGND VGND VPWR VPWR _08480_/B sky130_fd_sc_hd__nand2_1
X_10510_ _10512_/A _10510_/B VGND VGND VPWR VPWR _14431_/D sky130_fd_sc_hd__nor2_1
XFILLER_10_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11490_ _11490_/A VGND VGND VPWR VPWR _13831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10441_ _10441_/A _10460_/A VGND VGND VPWR VPWR _10449_/A sky130_fd_sc_hd__and2_1
XFILLER_137_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10372_ _10432_/A _10432_/B _10376_/C _10415_/A _10378_/B VGND VGND VPWR VPWR _14214_/D
+ sky130_fd_sc_hd__o221a_1
X_13160_ _13554_/CLK _13160_/D _12609_/A VGND VGND VPWR VPWR _13160_/Q sky130_fd_sc_hd__dfrtp_1
X_12111_ _14471_/Q _11972_/X _12117_/S VGND VGND VPWR VPWR _12112_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13091_ _13562_/CLK hold310/X VGND VGND VPWR VPWR _13091_/Q sky130_fd_sc_hd__dfxtp_1
X_12042_ _12076_/A VGND VGND VPWR VPWR _12093_/S sky130_fd_sc_hd__buf_2
XFILLER_123_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold290 hold290/A VGND VGND VPWR VPWR hold290/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_49_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13993_ _14707_/CLK _13993_/D VGND VGND VPWR VPWR _13993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12944_ _13280_/CLK _12944_/D VGND VGND VPWR VPWR hold258/A sky130_fd_sc_hd__dfxtp_1
XFILLER_92_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _14678_/CLK _12875_/D VGND VGND VPWR VPWR _12875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _14615_/CLK _14614_/D VGND VGND VPWR VPWR _14614_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _13583_/Q _11828_/B VGND VGND VPWR VPWR _11827_/A sky130_fd_sc_hd__and2_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _14652_/CLK _14545_/D VGND VGND VPWR VPWR _14545_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _11757_/A VGND VGND VPWR VPWR _14069_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_134_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _14210_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10708_ _10708_/A VGND VGND VPWR VPWR _12932_/D sky130_fd_sc_hd__clkbuf_1
X_14476_ _14543_/CLK _14476_/D VGND VGND VPWR VPWR _14476_/Q sky130_fd_sc_hd__dfxtp_1
X_11688_ _11688_/A VGND VGND VPWR VPWR _14026_/D sky130_fd_sc_hd__clkbuf_1
X_13427_ _14679_/CLK hold84/X VGND VGND VPWR VPWR _13427_/Q sky130_fd_sc_hd__dfxtp_2
X_10639_ _13962_/Q _13965_/Q _13936_/Q VGND VGND VPWR VPWR _10640_/B sky130_fd_sc_hd__o21ai_1
XFILLER_155_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13358_ _13434_/CLK _13358_/D repeater56/X VGND VGND VPWR VPWR _13358_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_127_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12309_ _14570_/Q _11991_/X _12313_/S VGND VGND VPWR VPWR _12310_/A sky130_fd_sc_hd__mux2_1
X_13289_ _13296_/CLK hold338/X VGND VGND VPWR VPWR _13289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07850_ _07858_/D _07850_/B VGND VGND VPWR VPWR _07850_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_68_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06801_ _06813_/A _06811_/A VGND VGND VPWR VPWR _06807_/A sky130_fd_sc_hd__xnor2_1
XFILLER_84_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07781_ _07766_/X _07780_/Y _07781_/S VGND VGND VPWR VPWR _07782_/A sky130_fd_sc_hd__mux2_1
Xinput3 data_i[11] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__buf_8
X_09520_ _09513_/A _09514_/X _09534_/B VGND VGND VPWR VPWR _09520_/Y sky130_fd_sc_hd__a21oi_1
X_06732_ _06895_/A VGND VGND VPWR VPWR _06871_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09451_ _13601_/Q _09451_/B VGND VGND VPWR VPWR _09452_/B sky130_fd_sc_hd__or2_1
X_06663_ _06656_/X _06661_/X _07909_/A VGND VGND VPWR VPWR _06664_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08402_ _13097_/Q _13378_/Q _08406_/S VGND VGND VPWR VPWR _08403_/A sky130_fd_sc_hd__mux2_1
X_06594_ _12897_/Q _06590_/A _06593_/Y _06542_/X VGND VGND VPWR VPWR _12897_/D sky130_fd_sc_hd__o211a_1
X_09382_ _09382_/A _09382_/B VGND VGND VPWR VPWR _09385_/A sky130_fd_sc_hd__nand2_1
XFILLER_101_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08333_ _08333_/A _08333_/B VGND VGND VPWR VPWR _13381_/D sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_125_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _13843_/CLK sky130_fd_sc_hd__clkbuf_16
X_08264_ _13367_/Q _08268_/B VGND VGND VPWR VPWR _08265_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07215_ _07215_/A _07215_/B VGND VGND VPWR VPWR _07215_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_137_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08195_ _08195_/A VGND VGND VPWR VPWR _13360_/D sky130_fd_sc_hd__clkbuf_1
X_07146_ _07171_/B _07146_/B VGND VGND VPWR VPWR _07147_/B sky130_fd_sc_hd__xnor2_2
XFILLER_161_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07077_ _07077_/A _07077_/B _07077_/C VGND VGND VPWR VPWR _07078_/B sky130_fd_sc_hd__or3_1
XFILLER_134_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06028_ _06353_/A _12030_/C VGND VGND VPWR VPWR _14590_/D sky130_fd_sc_hd__nand2_1
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07979_ _07987_/A _07986_/A _06976_/A VGND VGND VPWR VPWR _07979_/X sky130_fd_sc_hd__o21a_1
XFILLER_28_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09718_ _09718_/A _09736_/A VGND VGND VPWR VPWR _09718_/Y sky130_fd_sc_hd__nand2_1
X_10990_ _13321_/Q _10907_/X _10983_/X _10989_/Y VGND VGND VPWR VPWR _13321_/D sky130_fd_sc_hd__o22a_1
XFILLER_142_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09649_ _13420_/Q _13618_/Q _09653_/S VGND VGND VPWR VPWR _09650_/A sky130_fd_sc_hd__mux2_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _14737_/CLK hold488/X _12609_/A VGND VGND VPWR VPWR _12661_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11611_/A VGND VGND VPWR VPWR _13982_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12591_ _12616_/B _12591_/B _12591_/C _12591_/D VGND VGND VPWR VPWR _12591_/X sky130_fd_sc_hd__or4_1
XFILLER_24_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_116_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _13622_/CLK sky130_fd_sc_hd__clkbuf_16
X_14330_ _14696_/CLK hold432/X VGND VGND VPWR VPWR hold398/A sky130_fd_sc_hd__dfxtp_1
X_11542_ _11542_/A VGND VGND VPWR VPWR _13854_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14261_ _14707_/CLK _14261_/D VGND VGND VPWR VPWR _14261_/Q sky130_fd_sc_hd__dfxtp_1
X_11473_ _13826_/Q _11472_/X _11479_/S VGND VGND VPWR VPWR _11474_/A sky130_fd_sc_hd__mux2_1
X_13212_ _13702_/CLK _13212_/D VGND VGND VPWR VPWR _13212_/Q sky130_fd_sc_hd__dfxtp_1
X_10424_ _10374_/A _10431_/A _10423_/X _10416_/B VGND VGND VPWR VPWR _10426_/C sky130_fd_sc_hd__a31o_1
X_14192_ _14610_/CLK _14192_/D VGND VGND VPWR VPWR hold299/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13143_ _13535_/CLK _13143_/D repeater57/X VGND VGND VPWR VPWR _13143_/Q sky130_fd_sc_hd__dfrtp_1
X_10355_ _13780_/Q _13781_/Q VGND VGND VPWR VPWR _10359_/B sky130_fd_sc_hd__nor2_1
XFILLER_152_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _10285_/X _10282_/X _10286_/S VGND VGND VPWR VPWR _10287_/A sky130_fd_sc_hd__mux2_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _14636_/CLK hold494/X VGND VGND VPWR VPWR _13074_/Q sky130_fd_sc_hd__dfxtp_1
X_12025_ _12025_/A VGND VGND VPWR VPWR _12025_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13976_ _13978_/CLK _13976_/D VGND VGND VPWR VPWR _13976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12927_ _13263_/CLK _12927_/D VGND VGND VPWR VPWR hold226/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12858_ _13686_/CLK _12858_/D VGND VGND VPWR VPWR hold70/A sky130_fd_sc_hd__dfxtp_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11809_ _13575_/Q _11817_/B VGND VGND VPWR VPWR _11810_/A sky130_fd_sc_hd__and2_1
XFILLER_15_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_107_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _13621_/CLK sky130_fd_sc_hd__clkbuf_16
X_12789_ _13570_/CLK _12789_/D VGND VGND VPWR VPWR hold402/A sky130_fd_sc_hd__dfxtp_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14528_ _14557_/CLK _14528_/D VGND VGND VPWR VPWR _14528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14459_ _14615_/CLK _14459_/D VGND VGND VPWR VPWR _14459_/Q sky130_fd_sc_hd__dfxtp_1
X_07000_ _07001_/B _07001_/C _07001_/A VGND VGND VPWR VPWR _07000_/X sky130_fd_sc_hd__a21o_1
XFILLER_115_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08951_ _08951_/A _08951_/B _08951_/C VGND VGND VPWR VPWR _08952_/B sky130_fd_sc_hd__and3_1
XFILLER_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07902_ _13266_/Q _07902_/B VGND VGND VPWR VPWR _07903_/B sky130_fd_sc_hd__or2_1
X_08882_ _08895_/B _08895_/C VGND VGND VPWR VPWR _08883_/B sky130_fd_sc_hd__nor2_1
XFILLER_96_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07833_ _07833_/A _07833_/B _07828_/B VGND VGND VPWR VPWR _07858_/A sky130_fd_sc_hd__or3b_2
XFILLER_57_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07764_ _07764_/A _07764_/B _07764_/C VGND VGND VPWR VPWR _07765_/B sky130_fd_sc_hd__and3_1
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09503_ _13608_/Q _09530_/B VGND VGND VPWR VPWR _09509_/D sky130_fd_sc_hd__xnor2_1
X_06715_ _06703_/X _07832_/B _06714_/X VGND VGND VPWR VPWR _13002_/D sky130_fd_sc_hd__a21o_1
X_07695_ _07695_/A _07695_/B VGND VGND VPWR VPWR _07697_/A sky130_fd_sc_hd__xnor2_1
XFILLER_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09434_ _09454_/A _09454_/B _09454_/C VGND VGND VPWR VPWR _09443_/B sky130_fd_sc_hd__or3_1
XFILLER_25_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06646_ _13345_/Q _13343_/Q _06704_/S VGND VGND VPWR VPWR _06646_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09365_ _09365_/A _13589_/Q VGND VGND VPWR VPWR _09366_/B sky130_fd_sc_hd__nand2_1
X_06577_ _12892_/Q _12893_/Q VGND VGND VPWR VPWR _06584_/D sky130_fd_sc_hd__and2_1
X_08316_ _08316_/A _08316_/B VGND VGND VPWR VPWR _13376_/D sky130_fd_sc_hd__nor2_1
XANTENNA_30 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09296_ _09296_/A VGND VGND VPWR VPWR _12776_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_41 _13334_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 hold502/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 _13090_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08247_ _08247_/A _08247_/B VGND VGND VPWR VPWR _08247_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_74 _11092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_85 _13329_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_96 _13700_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08178_ _08261_/A _10310_/A _08116_/X _13427_/Q VGND VGND VPWR VPWR _08178_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_137_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07129_ _07151_/B _07128_/B _07128_/C VGND VGND VPWR VPWR _07130_/B sky130_fd_sc_hd__a21oi_1
XFILLER_133_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10140_ _10149_/B VGND VGND VPWR VPWR _14140_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10071_ _13919_/Q _10056_/X _10063_/A VGND VGND VPWR VPWR _14042_/D sky130_fd_sc_hd__a21o_1
XFILLER_102_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13830_ _14713_/CLK _13830_/D VGND VGND VPWR VPWR _13830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13761_ _14709_/CLK _13761_/D VGND VGND VPWR VPWR _13761_/Q sky130_fd_sc_hd__dfxtp_1
X_10973_ _14747_/Q VGND VGND VPWR VPWR _11190_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12712_ _13593_/CLK _12712_/D VGND VGND VPWR VPWR hold458/A sky130_fd_sc_hd__dfxtp_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13692_ _13855_/CLK _13692_/D repeater57/X VGND VGND VPWR VPWR _13692_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12643_ _12643_/A _12645_/B VGND VGND VPWR VPWR _12643_/X sky130_fd_sc_hd__or2_1
XFILLER_43_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12574_ _14740_/Q VGND VGND VPWR VPWR _12625_/A sky130_fd_sc_hd__inv_2
X_14313_ _14510_/CLK _14313_/D VGND VGND VPWR VPWR _14313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11525_ _13623_/Q _11529_/B VGND VGND VPWR VPWR _11526_/A sky130_fd_sc_hd__and2_1
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14244_ _14726_/CLK _14244_/D VGND VGND VPWR VPWR _14244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11456_ _14696_/Q VGND VGND VPWR VPWR _11456_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10407_ _10407_/A _10407_/B _10405_/Y VGND VGND VPWR VPWR _10411_/C sky130_fd_sc_hd__or3b_1
XFILLER_124_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14175_ _14209_/CLK _14175_/D VGND VGND VPWR VPWR _14175_/Q sky130_fd_sc_hd__dfxtp_1
X_11387_ _11387_/A VGND VGND VPWR VPWR _13786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13126_ _14645_/CLK _13708_/Q VGND VGND VPWR VPWR hold64/A sky130_fd_sc_hd__dfxtp_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10338_ _10339_/A hold131/A _10339_/C VGND VGND VPWR VPWR _10340_/A sky130_fd_sc_hd__o21a_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _13562_/CLK _13057_/D VGND VGND VPWR VPWR hold378/A sky130_fd_sc_hd__dfxtp_1
X_10269_ _10266_/X _14357_/D _10269_/S VGND VGND VPWR VPWR _10270_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12008_ _14312_/Q _12007_/X _12014_/S VGND VGND VPWR VPWR _12009_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13959_ _13963_/CLK _13959_/D VGND VGND VPWR VPWR _13959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06500_ _06500_/A _06500_/B VGND VGND VPWR VPWR _06500_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07480_ _13148_/Q _09228_/B VGND VGND VPWR VPWR _07493_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06431_ _12879_/Q _06450_/B VGND VGND VPWR VPWR _06433_/A sky130_fd_sc_hd__or2_1
X_06362_ _14643_/Q _12340_/B _14633_/D _14639_/Q VGND VGND VPWR VPWR _14428_/D sky130_fd_sc_hd__a22o_1
X_09150_ _09106_/X _09156_/B _09149_/Y _07396_/X VGND VGND VPWR VPWR _13533_/D sky130_fd_sc_hd__a31o_1
XFILLER_147_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08101_ _08164_/A VGND VGND VPWR VPWR _08199_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06293_ _14187_/Q _14179_/Q _10110_/A VGND VGND VPWR VPWR _06293_/X sky130_fd_sc_hd__mux2_1
X_09081_ _09081_/A VGND VGND VPWR VPWR _12773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08032_ _12954_/Q _13254_/Q _08040_/S VGND VGND VPWR VPWR _08033_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14751__62 VGND VGND VPWR VPWR _14751__62/HI data_o[25] sky130_fd_sc_hd__conb_1
XFILLER_131_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09983_ _09983_/A VGND VGND VPWR VPWR _13705_/D sky130_fd_sc_hd__clkbuf_1
X_08934_ _08959_/B _08934_/B VGND VGND VPWR VPWR _08935_/B sky130_fd_sc_hd__xnor2_1
XFILLER_69_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08865_ _08865_/A _08865_/B _08865_/C VGND VGND VPWR VPWR _08866_/B sky130_fd_sc_hd__or3_1
XFILLER_96_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07816_ _07815_/B _07815_/C _07815_/A VGND VGND VPWR VPWR _07816_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08796_ _08794_/Y _08795_/X _08735_/X VGND VGND VPWR VPWR _13466_/D sky130_fd_sc_hd__o21bai_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07747_ _07747_/A _07772_/D VGND VGND VPWR VPWR _07748_/B sky130_fd_sc_hd__nand2_1
XFILLER_41_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07678_ _07708_/A _07708_/B VGND VGND VPWR VPWR _07680_/A sky130_fd_sc_hd__xnor2_1
XFILLER_13_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09417_ _09408_/A _09417_/B _13595_/Q VGND VGND VPWR VPWR _09420_/B sky130_fd_sc_hd__and3b_1
X_06629_ _13036_/Q VGND VGND VPWR VPWR _06630_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09348_ _13310_/Q _13548_/Q _09354_/S VGND VGND VPWR VPWR _09349_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09279_ _09276_/Y _09277_/X _09272_/A _09273_/Y VGND VGND VPWR VPWR _09279_/X sky130_fd_sc_hd__a211o_1
XFILLER_154_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11310_ _14514_/Q VGND VGND VPWR VPWR _11310_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12290_ _12290_/A VGND VGND VPWR VPWR _14561_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11241_ _10944_/A _11238_/Y _11240_/Y _10929_/A VGND VGND VPWR VPWR _11242_/B sky130_fd_sc_hd__a211o_1
XFILLER_4_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11172_ _11172_/A _11155_/X VGND VGND VPWR VPWR _11172_/X sky130_fd_sc_hd__or2b_1
XFILLER_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10123_ _06145_/C _06146_/Y _10119_/S _10111_/X VGND VGND VPWR VPWR _14204_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10054_ _14038_/D _10062_/B VGND VGND VPWR VPWR _10060_/A sky130_fd_sc_hd__and2_1
XFILLER_0_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13813_ _13843_/CLK _13813_/D VGND VGND VPWR VPWR _13813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13744_ _13843_/CLK hold181/X VGND VGND VPWR VPWR _13843_/D sky130_fd_sc_hd__dfxtp_1
X_10956_ _14597_/Q _14559_/Q _14490_/Q _14442_/Q _11208_/A _11209_/A VGND VGND VPWR
+ VPWR _10957_/A sky130_fd_sc_hd__mux4_1
XFILLER_31_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13675_ _14251_/CLK _13675_/D repeater56/X VGND VGND VPWR VPWR _13675_/Q sky130_fd_sc_hd__dfrtp_1
X_10887_ _13160_/Q _10891_/B VGND VGND VPWR VPWR _10888_/A sky130_fd_sc_hd__and2_1
X_12626_ _14740_/Q _12626_/B VGND VGND VPWR VPWR _12626_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12557_ _12557_/A VGND VGND VPWR VPWR _14723_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11508_ _13837_/Q _11507_/X _11511_/S VGND VGND VPWR VPWR _11509_/A sky130_fd_sc_hd__mux2_1
X_12488_ _12496_/A _12496_/B input10/X VGND VGND VPWR VPWR _12489_/A sky130_fd_sc_hd__and3_1
Xhold108 hold108/A VGND VGND VPWR VPWR hold108/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14227_ _14737_/CLK _14227_/D VGND VGND VPWR VPWR _14227_/Q sky130_fd_sc_hd__dfxtp_1
Xhold119 hold119/A VGND VGND VPWR VPWR hold119/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_11439_ _11439_/A VGND VGND VPWR VPWR _13810_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14158_ _14159_/CLK hold272/X VGND VGND VPWR VPWR hold215/A sky130_fd_sc_hd__dfxtp_1
XFILLER_113_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13109_ _14636_/CLK _13109_/D VGND VGND VPWR VPWR _13109_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _06976_/X _06979_/Y _06897_/X VGND VGND VPWR VPWR _13025_/D sky130_fd_sc_hd__a21o_1
X_14089_ _14098_/CLK _14089_/D VGND VGND VPWR VPWR _14089_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05931_ _13740_/Q _13741_/Q _13742_/Q _13743_/Q VGND VGND VPWR VPWR _05934_/A sky130_fd_sc_hd__or4_1
XFILLER_67_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08650_ _13449_/Q _08650_/B VGND VGND VPWR VPWR _08651_/B sky130_fd_sc_hd__or2_1
XFILLER_67_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07601_ _07601_/A _07620_/A VGND VGND VPWR VPWR _07602_/B sky130_fd_sc_hd__or2_1
X_08581_ _08581_/A _08581_/B VGND VGND VPWR VPWR _08582_/C sky130_fd_sc_hd__and2_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07532_ _07532_/A _07532_/B _07532_/C _07530_/C VGND VGND VPWR VPWR _07533_/B sky130_fd_sc_hd__or4b_1
XFILLER_81_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07463_ _09207_/B VGND VGND VPWR VPWR _07513_/B sky130_fd_sc_hd__clkbuf_2
X_09202_ _09205_/A _09220_/B VGND VGND VPWR VPWR _09202_/X sky130_fd_sc_hd__or2_1
XFILLER_50_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06414_ _06410_/X _06554_/B _06427_/S VGND VGND VPWR VPWR _06513_/B sky130_fd_sc_hd__mux2_2
XFILLER_10_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07394_ _07414_/A _07394_/B VGND VGND VPWR VPWR _07394_/X sky130_fd_sc_hd__xor2_1
X_09133_ _09114_/A _09119_/Y _09120_/Y _09134_/C _09134_/D VGND VGND VPWR VPWR _09135_/B
+ sky130_fd_sc_hd__a2111o_1
X_06345_ _14109_/Q _14093_/Q _06345_/S VGND VGND VPWR VPWR _06346_/A sky130_fd_sc_hd__mux2_1
X_06276_ _06276_/A VGND VGND VPWR VPWR _13956_/D sky130_fd_sc_hd__clkbuf_1
X_09064_ _13230_/Q _13459_/Q _09064_/S VGND VGND VPWR VPWR _09065_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08015_ _13282_/Q _08015_/B VGND VGND VPWR VPWR _08016_/B sky130_fd_sc_hd__or2_1
XFILLER_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09966_ hold456/X _13695_/Q _09968_/S VGND VGND VPWR VPWR _09967_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08917_ _08939_/B _08916_/B _08916_/C VGND VGND VPWR VPWR _08918_/B sky130_fd_sc_hd__a21oi_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _13697_/Q _09893_/A _09893_/B _09672_/Y VGND VGND VPWR VPWR _09897_/X sky130_fd_sc_hd__a31o_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_96_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _13681_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08848_ _13519_/D VGND VGND VPWR VPWR _08929_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ _13464_/Q _09569_/B VGND VGND VPWR VPWR _08779_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10810_ _13025_/Q _10812_/B VGND VGND VPWR VPWR _10811_/A sky130_fd_sc_hd__and2_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _11790_/A VGND VGND VPWR VPWR _14088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10741_ _10741_/A VGND VGND VPWR VPWR _12947_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13460_ _13698_/CLK _13460_/D repeater57/X VGND VGND VPWR VPWR _13460_/Q sky130_fd_sc_hd__dfrtp_2
X_10672_ _14341_/Q _10671_/C _14342_/Q VGND VGND VPWR VPWR _10673_/C sky130_fd_sc_hd__a21o_1
XFILLER_139_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12411_ _12411_/A VGND VGND VPWR VPWR _14639_/D sky130_fd_sc_hd__clkbuf_1
X_13391_ _14012_/CLK hold223/X VGND VGND VPWR VPWR _13391_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_20_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _14082_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_126_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12342_ _12342_/A _12342_/B VGND VGND VPWR VPWR _12377_/A sky130_fd_sc_hd__nor2_4
XFILLER_5_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12273_ _12273_/A VGND VGND VPWR VPWR _14551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14012_ _14012_/CLK _14012_/D VGND VGND VPWR VPWR _14012_/Q sky130_fd_sc_hd__dfxtp_1
X_11224_ _11224_/A VGND VGND VPWR VPWR _12647_/A sky130_fd_sc_hd__buf_2
XFILLER_135_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11155_ _11155_/A VGND VGND VPWR VPWR _11155_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10106_ _10106_/A VGND VGND VPWR VPWR _14142_/D sky130_fd_sc_hd__inv_2
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11086_ _11224_/A VGND VGND VPWR VPWR _11086_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_87_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _13520_/CLK sky130_fd_sc_hd__clkbuf_16
X_10037_ _06075_/D _06259_/Y _13965_/D _10029_/X VGND VGND VPWR VPWR _13973_/D sky130_fd_sc_hd__a22o_1
XFILLER_76_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11988_ _14516_/Q VGND VGND VPWR VPWR _11988_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13727_ _13727_/CLK hold313/X VGND VGND VPWR VPWR _13727_/Q sky130_fd_sc_hd__dfxtp_1
X_10939_ _11155_/A VGND VGND VPWR VPWR _10944_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13658_ _14679_/CLK _13658_/D VGND VGND VPWR VPWR _13658_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12609_ _12609_/A VGND VGND VPWR VPWR _12609_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13589_ _14010_/CLK _13589_/D repeater56/X VGND VGND VPWR VPWR _13589_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_11_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _13027_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06130_ _14204_/Q _14202_/Q _10107_/A VGND VGND VPWR VPWR _06130_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06061_ _06060_/X _06056_/X _10019_/A VGND VGND VPWR VPWR _06062_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09820_ _13680_/Q _09821_/B VGND VGND VPWR VPWR _09822_/A sky130_fd_sc_hd__and2_1
XFILLER_141_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09751_ _13672_/Q _09739_/B _09750_/X VGND VGND VPWR VPWR _09751_/Y sky130_fd_sc_hd__o21ai_1
X_06963_ _13022_/Q _08020_/B _06968_/A _06967_/A VGND VGND VPWR VPWR _06964_/B sky130_fd_sc_hd__a22o_1
XFILLER_67_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_78_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _14679_/CLK sky130_fd_sc_hd__clkbuf_16
X_08702_ _08709_/A _08702_/B VGND VGND VPWR VPWR _08714_/C sky130_fd_sc_hd__nand2_1
XFILLER_100_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05914_ _10050_/S VGND VGND VPWR VPWR _13935_/D sky130_fd_sc_hd__buf_2
X_09682_ _09682_/A _09682_/B VGND VGND VPWR VPWR _09683_/B sky130_fd_sc_hd__xnor2_1
X_06894_ _08008_/B VGND VGND VPWR VPWR _06895_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_39_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08633_ _08633_/A VGND VGND VPWR VPWR _08633_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _08578_/A _08564_/B VGND VGND VPWR VPWR _08581_/A sky130_fd_sc_hd__or2_1
XFILLER_35_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07515_ _07515_/A _07515_/B VGND VGND VPWR VPWR _07532_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08495_ _13438_/Q _08495_/B VGND VGND VPWR VPWR _08512_/A sky130_fd_sc_hd__nor2_1
XFILLER_50_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07446_ _07411_/X _07441_/Y _07454_/B _07445_/X VGND VGND VPWR VPWR _13145_/D sky130_fd_sc_hd__a31o_1
XFILLER_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07377_ _07350_/A _07375_/B _07364_/B _07374_/B VGND VGND VPWR VPWR _09139_/C sky130_fd_sc_hd__a31o_1
XFILLER_108_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09116_ _09120_/B _09115_/Y _09116_/S VGND VGND VPWR VPWR _09117_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06328_ _14379_/Q _14423_/D VGND VGND VPWR VPWR _06328_/X sky130_fd_sc_hd__and2_1
XFILLER_163_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09047_ _13223_/Q _13452_/Q _09051_/S VGND VGND VPWR VPWR _09048_/A sky130_fd_sc_hd__mux2_1
X_06259_ _06259_/A _06259_/B VGND VGND VPWR VPWR _06259_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold450 data_i[3] VGND VGND VPWR VPWR input20/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold461 hold461/A VGND VGND VPWR VPWR hold461/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_145_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold472 hold472/A VGND VGND VPWR VPWR hold472/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold483 hold483/A VGND VGND VPWR VPWR hold483/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_78_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold494 hold494/A VGND VGND VPWR VPWR hold494/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09949_ _13498_/Q _13687_/Q _09957_/S VGND VGND VPWR VPWR _09950_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_69_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _13555_/CLK sky130_fd_sc_hd__clkbuf_16
X_12960_ _13263_/CLK hold226/X VGND VGND VPWR VPWR _12960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11911_ _11911_/A VGND VGND VPWR VPWR _14262_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12891_ _12970_/CLK _12891_/D hold1/X VGND VGND VPWR VPWR _12891_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _14644_/CLK hold136/X VGND VGND VPWR VPWR _14630_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _12150_/A _12095_/B VGND VGND VPWR VPWR _11877_/A sky130_fd_sc_hd__nor2_8
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _14652_/CLK _14561_/D VGND VGND VPWR VPWR _14561_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11773_ _11773_/A VGND VGND VPWR VPWR _14081_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _14010_/CLK _13512_/D VGND VGND VPWR VPWR _13710_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_14_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10724_ _10724_/A VGND VGND VPWR VPWR _12939_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _14492_/CLK _14492_/D VGND VGND VPWR VPWR _14492_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13443_ _13702_/CLK _13443_/D repeater56/X VGND VGND VPWR VPWR _13443_/Q sky130_fd_sc_hd__dfrtp_1
X_10655_ _14320_/Q _14327_/Q VGND VGND VPWR VPWR _10673_/B sky130_fd_sc_hd__nor2_1
XFILLER_155_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13374_ _13377_/CLK _13374_/D repeater57/X VGND VGND VPWR VPWR _13374_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10586_ _13386_/Q _13434_/Q _13387_/Q _07343_/X VGND VGND VPWR VPWR _13386_/D sky130_fd_sc_hd__o31a_1
XFILLER_139_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12325_ _12325_/A VGND VGND VPWR VPWR _14577_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12256_ _12256_/A VGND VGND VPWR VPWR _14543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11207_ _11207_/A VGND VGND VPWR VPWR _11207_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12187_ _12187_/A VGND VGND VPWR VPWR _14504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11138_ _11209_/A VGND VGND VPWR VPWR _11138_/X sky130_fd_sc_hd__buf_4
XFILLER_122_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11069_ _14022_/Q _13988_/Q _13828_/Q _14540_/Q _11010_/X _11011_/X VGND VGND VPWR
+ VPWR _11070_/A sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_0_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _14510_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07300_ _07224_/A _07298_/X _07299_/X _07227_/X _07372_/S _07327_/A VGND VGND VPWR
+ VPWR _07311_/B sky130_fd_sc_hd__mux4_1
X_08280_ _13369_/Q _08281_/B VGND VGND VPWR VPWR _08282_/A sky130_fd_sc_hd__and2_1
X_07231_ _13167_/Q _07327_/A VGND VGND VPWR VPWR _07231_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07162_ _07163_/A _07203_/C _07163_/C VGND VGND VPWR VPWR _07164_/A sky130_fd_sc_hd__a21oi_1
XFILLER_118_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06113_ _13937_/D _13938_/D _13939_/D _13940_/D VGND VGND VPWR VPWR _06114_/C sky130_fd_sc_hd__or4_1
X_07093_ _07093_/A _07093_/B _07093_/C VGND VGND VPWR VPWR _07107_/C sky130_fd_sc_hd__nor3_2
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06044_ _10601_/A _06044_/B VGND VGND VPWR VPWR _12400_/C sky130_fd_sc_hd__nor2_1
XFILLER_160_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09803_ _09803_/A _09815_/A VGND VGND VPWR VPWR _09806_/A sky130_fd_sc_hd__or2b_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07995_ _07995_/A _07995_/B VGND VGND VPWR VPWR _07996_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09734_ _09735_/A _09819_/B _09736_/A VGND VGND VPWR VPWR _09734_/X sky130_fd_sc_hd__a21o_1
X_06946_ _13021_/Q _06954_/A VGND VGND VPWR VPWR _06950_/B sky130_fd_sc_hd__xor2_1
XFILLER_27_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09665_ _13710_/Q VGND VGND VPWR VPWR _09718_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06877_ _06877_/A _06877_/B VGND VGND VPWR VPWR _06877_/Y sky130_fd_sc_hd__nand2_1
XFILLER_131_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08616_ _08464_/X _08614_/Y _08615_/X VGND VGND VPWR VPWR _13446_/D sky130_fd_sc_hd__a21o_1
XFILLER_43_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _13396_/Q _13594_/Q _09598_/S VGND VGND VPWR VPWR _09597_/A sky130_fd_sc_hd__mux2_2
XFILLER_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _08645_/A _08545_/X _08546_/Y VGND VGND VPWR VPWR _08657_/B sky130_fd_sc_hd__o21ba_1
XFILLER_70_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08478_ _08478_/A VGND VGND VPWR VPWR _09383_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07429_ _07329_/Y _07428_/Y _07327_/X VGND VGND VPWR VPWR _07435_/B sky130_fd_sc_hd__o21ai_2
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10440_ hold79/A VGND VGND VPWR VPWR _10460_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_137_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10371_ _10432_/A _10386_/A _10374_/A VGND VGND VPWR VPWR _10378_/B sky130_fd_sc_hd__nand3_1
XFILLER_108_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12110_ _12110_/A VGND VGND VPWR VPWR _14470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13090_ _13562_/CLK hold378/X VGND VGND VPWR VPWR _13090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12041_ _12621_/A _12619_/A _12041_/C VGND VGND VPWR VPWR _12076_/A sky130_fd_sc_hd__nand3b_4
XFILLER_105_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold280 hold280/A VGND VGND VPWR VPWR hold280/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_151_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold291 hold291/A VGND VGND VPWR VPWR hold291/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13992_ _14707_/CLK _13992_/D VGND VGND VPWR VPWR _13992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ _13280_/CLK _12943_/D VGND VGND VPWR VPWR hold255/A sky130_fd_sc_hd__dfxtp_1
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ _14688_/CLK _12874_/D VGND VGND VPWR VPWR _12874_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ _14615_/CLK _14613_/D VGND VGND VPWR VPWR _14613_/Q sky130_fd_sc_hd__dfxtp_1
X_11825_ _11825_/A VGND VGND VPWR VPWR _14104_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _14707_/CLK _14544_/D VGND VGND VPWR VPWR _14544_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11756_ _11348_/X _14069_/Q _11758_/S VGND VGND VPWR VPWR _11757_/A sky130_fd_sc_hd__mux2_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _12889_/Q _10709_/B VGND VGND VPWR VPWR _10708_/A sky130_fd_sc_hd__and2_1
X_14475_ _14602_/CLK _14475_/D VGND VGND VPWR VPWR _14475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11687_ _14026_/Q _11491_/X _11689_/S VGND VGND VPWR VPWR _11688_/A sky130_fd_sc_hd__mux2_1
X_13426_ _13657_/CLK hold206/X VGND VGND VPWR VPWR _13426_/Q sky130_fd_sc_hd__dfxtp_1
X_10638_ _13962_/Q _13965_/Q VGND VGND VPWR VPWR _13913_/D sky130_fd_sc_hd__xor2_1
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13357_ _13657_/CLK _13357_/D hold1/X VGND VGND VPWR VPWR _13357_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10569_ _10570_/A _10570_/B _10570_/C VGND VGND VPWR VPWR _10575_/B sky130_fd_sc_hd__a21o_1
XFILLER_143_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12308_ _12308_/A VGND VGND VPWR VPWR _14569_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13288_ _13525_/CLK hold58/X VGND VGND VPWR VPWR _13288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12239_ _12261_/A VGND VGND VPWR VPWR _12248_/S sky130_fd_sc_hd__buf_2
XFILLER_111_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06800_ _06800_/A _06800_/B VGND VGND VPWR VPWR _06811_/A sky130_fd_sc_hd__nor2_1
XFILLER_111_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07780_ _07791_/A _07780_/B VGND VGND VPWR VPWR _07780_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_83_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput4 data_i[12] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06731_ _06731_/A _06731_/B VGND VGND VPWR VPWR _06731_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09450_ _13601_/Q _09450_/B VGND VGND VPWR VPWR _09460_/A sky130_fd_sc_hd__nand2_1
XFILLER_52_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06662_ _13032_/Q VGND VGND VPWR VPWR _07909_/A sky130_fd_sc_hd__buf_4
XFILLER_92_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08401_ _08401_/A VGND VGND VPWR VPWR _12732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09381_ _13592_/Q _09388_/B VGND VGND VPWR VPWR _09382_/B sky130_fd_sc_hd__nand2_1
X_06593_ _06593_/A VGND VGND VPWR VPWR _06593_/Y sky130_fd_sc_hd__inv_2
X_08332_ _08331_/A _08331_/B _08298_/X VGND VGND VPWR VPWR _08333_/B sky130_fd_sc_hd__o21ai_1
X_08263_ _13367_/Q _08268_/B VGND VGND VPWR VPWR _08265_/A sky130_fd_sc_hd__and2_1
XFILLER_137_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07214_ _07214_/A _07214_/B VGND VGND VPWR VPWR _07215_/B sky130_fd_sc_hd__xnor2_1
XFILLER_146_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08194_ _08188_/B _08193_/X _08215_/S VGND VGND VPWR VPWR _08195_/A sky130_fd_sc_hd__mux2_1
X_07145_ _07111_/A _07113_/B _07111_/B VGND VGND VPWR VPWR _07146_/B sky130_fd_sc_hd__o21ba_1
XFILLER_3_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07076_ _07077_/A _07077_/B _07077_/C VGND VGND VPWR VPWR _07101_/A sky130_fd_sc_hd__o21ai_2
XFILLER_160_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06027_ _14684_/Q _14686_/Q _06027_/C VGND VGND VPWR VPWR _12030_/C sky130_fd_sc_hd__or3_1
XFILLER_59_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07978_ _07987_/A _07986_/A VGND VGND VPWR VPWR _07978_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09717_ _14216_/Q _14214_/Q _09731_/A VGND VGND VPWR VPWR _09717_/X sky130_fd_sc_hd__mux2_1
X_06929_ _06951_/A _06928_/B _06836_/X VGND VGND VPWR VPWR _06929_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09648_ _09648_/A VGND VGND VPWR VPWR _12836_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _09579_/A _09579_/B _09579_/C VGND VGND VPWR VPWR _09579_/Y sky130_fd_sc_hd__nand3_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _13982_/Q _11459_/X _11612_/S VGND VGND VPWR VPWR _11611_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _12590_/A _14732_/Q VGND VGND VPWR VPWR _12591_/D sky130_fd_sc_hd__xor2_1
XFILLER_70_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11541_ _13630_/Q _11541_/B VGND VGND VPWR VPWR _11542_/A sky130_fd_sc_hd__and2_1
XFILLER_11_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14260_ _14707_/CLK _14260_/D VGND VGND VPWR VPWR _14260_/Q sky130_fd_sc_hd__dfxtp_1
X_11472_ _14701_/Q VGND VGND VPWR VPWR _11472_/X sky130_fd_sc_hd__buf_2
XFILLER_137_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13211_ _13596_/CLK hold437/X VGND VGND VPWR VPWR _13211_/Q sky130_fd_sc_hd__dfxtp_1
X_10423_ _10423_/A _10429_/C VGND VGND VPWR VPWR _10423_/X sky130_fd_sc_hd__or2_1
XFILLER_109_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14191_ _14693_/CLK _14191_/D VGND VGND VPWR VPWR _14191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13142_ _13532_/CLK _13142_/D repeater57/X VGND VGND VPWR VPWR _13142_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10354_ _13109_/D _13121_/D _10353_/X VGND VGND VPWR VPWR _13034_/D sky130_fd_sc_hd__o21a_1
XFILLER_2_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13073_ _13524_/CLK hold180/X VGND VGND VPWR VPWR _13073_/Q sky130_fd_sc_hd__dfxtp_1
X_10285_ _12874_/Q _14325_/Q _10593_/A VGND VGND VPWR VPWR _10285_/X sky130_fd_sc_hd__mux2_1
X_12024_ _12024_/A VGND VGND VPWR VPWR _14317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13975_ _14179_/CLK _13975_/D VGND VGND VPWR VPWR _13975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12926_ _12930_/CLK _12926_/D VGND VGND VPWR VPWR hold91/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12857_ _13805_/CLK _12857_/D VGND VGND VPWR VPWR hold303/A sky130_fd_sc_hd__dfxtp_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11808_ _11819_/A VGND VGND VPWR VPWR _11817_/B sky130_fd_sc_hd__clkbuf_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _13303_/CLK _12788_/D VGND VGND VPWR VPWR hold165/A sky130_fd_sc_hd__dfxtp_1
XFILLER_159_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11739_ _11313_/X _14061_/Q _11747_/S VGND VGND VPWR VPWR _11740_/A sky130_fd_sc_hd__mux2_1
X_14527_ _14555_/CLK _14527_/D VGND VGND VPWR VPWR _14527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14458_ _14615_/CLK _14458_/D VGND VGND VPWR VPWR _14458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13409_ _13617_/CLK hold495/X VGND VGND VPWR VPWR _13409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14389_ _14413_/CLK _14389_/D VGND VGND VPWR VPWR _14389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08950_ _08951_/A _08991_/C _08951_/C VGND VGND VPWR VPWR _08952_/A sky130_fd_sc_hd__a21oi_1
XFILLER_88_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07901_ _13266_/Q _07902_/B VGND VGND VPWR VPWR _07914_/A sky130_fd_sc_hd__nand2_1
X_08881_ _08881_/A _08881_/B _08881_/C VGND VGND VPWR VPWR _08895_/C sky130_fd_sc_hd__nor3_2
XFILLER_96_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07832_ _13256_/Q _07832_/B VGND VGND VPWR VPWR _07835_/A sky130_fd_sc_hd__nand2_2
XFILLER_38_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07763_ _07764_/A _07764_/B _07764_/C VGND VGND VPWR VPWR _07765_/A sky130_fd_sc_hd__a21oi_1
XFILLER_38_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09502_ _09502_/A VGND VGND VPWR VPWR _09502_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06714_ _07802_/A _06730_/B _06714_/C VGND VGND VPWR VPWR _06714_/X sky130_fd_sc_hd__and3_1
X_07694_ _13246_/D _13113_/Q VGND VGND VPWR VPWR _07695_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09433_ _09421_/A _09421_/B _09446_/C VGND VGND VPWR VPWR _09454_/C sky130_fd_sc_hd__o21a_1
XFILLER_64_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06645_ _13349_/Q _13347_/Q _06704_/S VGND VGND VPWR VPWR _06645_/X sky130_fd_sc_hd__mux2_1
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09364_ _09364_/A VGND VGND VPWR VPWR _12807_/D sky130_fd_sc_hd__clkbuf_1
X_06576_ _12892_/Q _06574_/X _06575_/Y VGND VGND VPWR VPWR _12892_/D sky130_fd_sc_hd__o21a_1
X_08315_ _13376_/Q _08312_/A _08338_/A VGND VGND VPWR VPWR _08316_/B sky130_fd_sc_hd__o21ai_1
XANTENNA_20 input26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09295_ _13286_/Q _13524_/Q _09299_/S VGND VGND VPWR VPWR _09296_/A sky130_fd_sc_hd__mux2_1
XANTENNA_31 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 _13319_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 input7/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08246_ _08236_/A _08245_/Y _08236_/B _08233_/A VGND VGND VPWR VPWR _08247_/B sky130_fd_sc_hd__a31o_1
XANTENNA_64 hold62/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_75 _11179_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_86 input4/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_97 _13700_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08177_ _08177_/A VGND VGND VPWR VPWR _10310_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07128_ _07151_/B _07128_/B _07128_/C VGND VGND VPWR VPWR _07153_/A sky130_fd_sc_hd__and3_1
XFILLER_107_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07059_ _07059_/A _07059_/B _07074_/B VGND VGND VPWR VPWR _07072_/A sky130_fd_sc_hd__or3_1
XFILLER_121_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10070_ _10070_/A VGND VGND VPWR VPWR _14044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13760_ _14710_/CLK _13760_/D VGND VGND VPWR VPWR _13760_/Q sky130_fd_sc_hd__dfxtp_1
X_10972_ _10972_/A VGND VGND VPWR VPWR _10972_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12711_ _13593_/CLK _12711_/D VGND VGND VPWR VPWR hold399/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13691_ _13855_/CLK _13691_/D repeater57/X VGND VGND VPWR VPWR _13691_/Q sky130_fd_sc_hd__dfrtp_2
X_12642_ _12642_/A VGND VGND VPWR VPWR _14745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12573_ _14741_/Q VGND VGND VPWR VPWR _12573_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14312_ _14510_/CLK _14312_/D VGND VGND VPWR VPWR _14312_/Q sky130_fd_sc_hd__dfxtp_1
X_11524_ _11524_/A VGND VGND VPWR VPWR _13842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14243_ _14726_/CLK _14243_/D VGND VGND VPWR VPWR _14243_/Q sky130_fd_sc_hd__dfxtp_1
X_11455_ _11455_/A VGND VGND VPWR VPWR _13820_/D sky130_fd_sc_hd__clkbuf_1
X_10406_ _10407_/A _10407_/B _10405_/Y VGND VGND VPWR VPWR _10421_/A sky130_fd_sc_hd__o21ba_1
X_14174_ _14201_/CLK _14174_/D VGND VGND VPWR VPWR _14174_/Q sky130_fd_sc_hd__dfxtp_1
X_11386_ _13717_/Q _11394_/B VGND VGND VPWR VPWR _11387_/A sky130_fd_sc_hd__and2_1
X_13125_ _14645_/CLK _13707_/Q VGND VGND VPWR VPWR hold79/A sky130_fd_sc_hd__dfxtp_2
XFILLER_125_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10337_ _14622_/Q _10337_/B VGND VGND VPWR VPWR _10339_/C sky130_fd_sc_hd__xnor2_1
XFILLER_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _13562_/CLK _13056_/D VGND VGND VPWR VPWR hold108/A sky130_fd_sc_hd__dfxtp_1
X_10268_ _10268_/A VGND VGND VPWR VPWR _14355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12007_ _12007_/A VGND VGND VPWR VPWR _12007_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_79_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10199_ _10208_/S VGND VGND VPWR VPWR _10206_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_93_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13958_ _13963_/CLK _13958_/D VGND VGND VPWR VPWR _13958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12909_ _14432_/CLK hold72/X VGND VGND VPWR VPWR _13031_/D sky130_fd_sc_hd__dfxtp_4
X_13889_ _14693_/CLK hold481/X VGND VGND VPWR VPWR _13889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06430_ _10346_/A _06446_/A _06524_/C _06429_/X VGND VGND VPWR VPWR _06450_/B sky130_fd_sc_hd__a31o_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06361_ _06361_/A VGND VGND VPWR VPWR _12340_/B sky130_fd_sc_hd__clkbuf_1
X_08100_ _13427_/Q VGND VGND VPWR VPWR _08164_/A sky130_fd_sc_hd__inv_2
X_09080_ _13237_/Q _13466_/Q _09587_/S VGND VGND VPWR VPWR _09081_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06292_ _06292_/A _06292_/B VGND VGND VPWR VPWR _06292_/Y sky130_fd_sc_hd__nand2_1
X_08031_ _10803_/A VGND VGND VPWR VPWR _08040_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09982_ _09977_/X _12404_/B _10596_/B VGND VGND VPWR VPWR _09983_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08933_ _08899_/A _08901_/B _08899_/B VGND VGND VPWR VPWR _08934_/B sky130_fd_sc_hd__o21ba_1
XFILLER_130_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08864_ _08865_/A _08865_/B _08865_/C VGND VGND VPWR VPWR _08889_/A sky130_fd_sc_hd__o21ai_2
XFILLER_57_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07815_ _07815_/A _07815_/B _07815_/C VGND VGND VPWR VPWR _07815_/Y sky130_fd_sc_hd__nand3_1
X_08795_ _08789_/A _08790_/X _08793_/Y _08733_/X VGND VGND VPWR VPWR _08795_/X sky130_fd_sc_hd__a31o_1
XFILLER_57_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07746_ _07746_/A _07746_/B VGND VGND VPWR VPWR _07748_/A sky130_fd_sc_hd__nor2_1
XFILLER_26_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07677_ _07689_/A _07677_/B VGND VGND VPWR VPWR _07708_/B sky130_fd_sc_hd__xnor2_1
XFILLER_25_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09416_ _09447_/A _09447_/B VGND VGND VPWR VPWR _09421_/A sky130_fd_sc_hd__or2_1
X_06628_ _07209_/A VGND VGND VPWR VPWR _13036_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_25_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09347_ _09347_/A VGND VGND VPWR VPWR _12799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06559_ _06537_/A _06548_/Y _06537_/B _06550_/A _06558_/X VGND VGND VPWR VPWR _06560_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_139_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09278_ _09272_/A _09273_/Y _09276_/Y _09277_/X VGND VGND VPWR VPWR _09278_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_21_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08229_ _08231_/B _08250_/C VGND VGND VPWR VPWR _08232_/B sky130_fd_sc_hd__and2_1
XFILLER_154_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11240_ _11240_/A _11240_/B VGND VGND VPWR VPWR _11240_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11171_ _14029_/Q _13995_/Q _13835_/Q _14547_/Q _11152_/X _11153_/X VGND VGND VPWR
+ VPWR _11172_/A sky130_fd_sc_hd__mux4_1
XFILLER_122_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10122_ _10122_/A VGND VGND VPWR VPWR _14203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10053_ _10062_/B VGND VGND VPWR VPWR _13908_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13812_ _13843_/CLK _13812_/D VGND VGND VPWR VPWR _13812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10955_ _12649_/B VGND VGND VPWR VPWR _10962_/A sky130_fd_sc_hd__buf_2
XFILLER_16_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13743_ _13843_/CLK hold155/X VGND VGND VPWR VPWR _13743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10886_ _10886_/A VGND VGND VPWR VPWR _13201_/D sky130_fd_sc_hd__clkbuf_1
X_13674_ _13680_/CLK _13674_/D repeater56/X VGND VGND VPWR VPWR _13674_/Q sky130_fd_sc_hd__dfrtp_1
X_12625_ _12625_/A _12625_/B VGND VGND VPWR VPWR _12631_/C sky130_fd_sc_hd__nor2_1
XFILLER_8_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12556_ _11359_/X _14723_/Q _12562_/S VGND VGND VPWR VPWR _12557_/A sky130_fd_sc_hd__mux2_1
X_11507_ _12010_/A VGND VGND VPWR VPWR _11507_/X sky130_fd_sc_hd__clkbuf_2
X_12487_ input29/X VGND VGND VPWR VPWR _12496_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_156_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold109 hold109/A VGND VGND VPWR VPWR hold109/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14226_ _14737_/CLK _14226_/D VGND VGND VPWR VPWR _14226_/Q sky130_fd_sc_hd__dfxtp_1
X_11438_ _13741_/Q _11438_/B VGND VGND VPWR VPWR _11439_/A sky130_fd_sc_hd__and2_1
XFILLER_160_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14157_ _14159_/CLK hold215/X VGND VGND VPWR VPWR _14157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11369_ _13894_/Q _11362_/X _11368_/Y VGND VGND VPWR VPWR _12022_/A sky130_fd_sc_hd__o21a_4
XFILLER_99_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13108_ _14636_/CLK _13108_/D VGND VGND VPWR VPWR _13108_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14088_ _14098_/CLK _14088_/D VGND VGND VPWR VPWR _14088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05930_ _13843_/D _13713_/Q _13714_/Q _13715_/Q VGND VGND VPWR VPWR _05935_/B sky130_fd_sc_hd__or4_1
X_13039_ _13039_/CLK _13039_/D VGND VGND VPWR VPWR _13039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07600_ _07613_/A _07622_/A _07627_/C VGND VGND VPWR VPWR _07620_/A sky130_fd_sc_hd__and3_1
XFILLER_26_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08580_ _08657_/A _08579_/X _08566_/B VGND VGND VPWR VPWR _08581_/B sky130_fd_sc_hd__o21a_1
XFILLER_82_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07531_ _07495_/X _07529_/Y _07530_/X _07499_/X VGND VGND VPWR VPWR _13154_/D sky130_fd_sc_hd__a31o_1
X_07462_ _07481_/A VGND VGND VPWR VPWR _09207_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09201_ _09210_/A _09201_/B VGND VGND VPWR VPWR _09220_/B sky130_fd_sc_hd__nand2_1
X_06413_ _13107_/D VGND VGND VPWR VPWR _06427_/S sky130_fd_sc_hd__inv_2
X_07393_ _07369_/X _07415_/B _07415_/A VGND VGND VPWR VPWR _07394_/B sky130_fd_sc_hd__a21o_1
X_09132_ _13530_/Q _09126_/B _09131_/X VGND VGND VPWR VPWR _09135_/A sky130_fd_sc_hd__a21oi_1
X_06344_ _06344_/A VGND VGND VPWR VPWR _14407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09063_ _09063_/A VGND VGND VPWR VPWR _12765_/D sky130_fd_sc_hd__clkbuf_1
X_06275_ _13810_/Q _13794_/Q _06281_/S VGND VGND VPWR VPWR _06276_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08014_ _13282_/Q _08015_/B VGND VGND VPWR VPWR _08016_/A sky130_fd_sc_hd__nand2_1
XFILLER_151_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09965_ _09965_/A VGND VGND VPWR VPWR _12868_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08916_ _08939_/B _08916_/B _08916_/C VGND VGND VPWR VPWR _08941_/A sky130_fd_sc_hd__and3_1
XFILLER_76_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _13697_/Q VGND VGND VPWR VPWR _09896_/Y sky130_fd_sc_hd__inv_2
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08847_ _08847_/A _08847_/B _08862_/B VGND VGND VPWR VPWR _08860_/A sky130_fd_sc_hd__or3_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08778_ _08776_/Y _08777_/X _08735_/X VGND VGND VPWR VPWR _13463_/D sky130_fd_sc_hd__o21bai_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07729_ _07729_/A _07729_/B VGND VGND VPWR VPWR _07731_/A sky130_fd_sc_hd__xor2_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10740_ _12904_/Q _10742_/B VGND VGND VPWR VPWR _10741_/A sky130_fd_sc_hd__and2_1
XFILLER_159_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10671_ _14341_/Q _14342_/Q _10671_/C VGND VGND VPWR VPWR _10671_/X sky130_fd_sc_hd__and3_1
X_12410_ _12418_/A _12418_/B input25/X VGND VGND VPWR VPWR _12411_/A sky130_fd_sc_hd__and3_1
XFILLER_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13390_ _13657_/CLK _13390_/D VGND VGND VPWR VPWR _13390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12341_ _12341_/A VGND VGND VPWR VPWR _14594_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12272_ _11359_/X _14551_/Q _12278_/S VGND VGND VPWR VPWR _12273_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14011_ _14012_/CLK _14011_/D VGND VGND VPWR VPWR _14011_/Q sky130_fd_sc_hd__dfxtp_1
X_11223_ _11223_/A _10960_/A VGND VGND VPWR VPWR _11223_/X sky130_fd_sc_hd__or2b_1
XFILLER_122_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11154_ _14028_/Q _13994_/Q _13834_/Q _14546_/Q _11152_/X _11153_/X VGND VGND VPWR
+ VPWR _11156_/A sky130_fd_sc_hd__mux4_1
XFILLER_1_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10105_ _10143_/A VGND VGND VPWR VPWR _14282_/D sky130_fd_sc_hd__inv_2
X_11085_ _11085_/A _11084_/X VGND VGND VPWR VPWR _11085_/X sky130_fd_sc_hd__or2b_1
XFILLER_103_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10036_ _06075_/C _06076_/Y _10032_/S _10024_/X VGND VGND VPWR VPWR _13972_/D sky130_fd_sc_hd__o22a_1
XFILLER_76_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11987_ _11987_/A VGND VGND VPWR VPWR _14305_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13726_ _13727_/CLK hold314/X VGND VGND VPWR VPWR _13726_/Q sky130_fd_sc_hd__dfxtp_1
X_10938_ _10938_/A VGND VGND VPWR VPWR _10938_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10869_ _10869_/A VGND VGND VPWR VPWR _13193_/D sky130_fd_sc_hd__clkbuf_1
X_13657_ _13657_/CLK _13657_/D VGND VGND VPWR VPWR _13657_/Q sky130_fd_sc_hd__dfxtp_1
X_12608_ _14733_/Q _12608_/B VGND VGND VPWR VPWR _12611_/A sky130_fd_sc_hd__and2_1
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13588_ _14530_/CLK hold476/X VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__dfxtp_1
XFILLER_129_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12539_ _11320_/X _14715_/Q _12543_/S VGND VGND VPWR VPWR _12540_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06060_ _13972_/Q _13970_/Q _10020_/A VGND VGND VPWR VPWR _06060_/X sky130_fd_sc_hd__mux2_1
X_14209_ _14209_/CLK _14209_/D VGND VGND VPWR VPWR _14209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06962_ _08015_/B VGND VGND VPWR VPWR _08020_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_98_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09750_ _13671_/Q _09722_/B _09739_/B _13672_/Q VGND VGND VPWR VPWR _09750_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05913_ _06273_/S VGND VGND VPWR VPWR _10050_/S sky130_fd_sc_hd__clkbuf_2
X_08701_ _13453_/Q _09511_/B VGND VGND VPWR VPWR _08702_/B sky130_fd_sc_hd__or2_1
X_09681_ _09681_/A _09680_/X VGND VGND VPWR VPWR _09682_/B sky130_fd_sc_hd__or2b_1
X_06893_ _08001_/B VGND VGND VPWR VPWR _08008_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08632_ _08617_/X _08629_/X _08630_/Y _08631_/X VGND VGND VPWR VPWR _13447_/D sky130_fd_sc_hd__a31o_1
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08563_ _08563_/A VGND VGND VPWR VPWR _13442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07514_ _13152_/Q _09212_/B VGND VGND VPWR VPWR _07515_/B sky130_fd_sc_hd__or2_1
XFILLER_63_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08494_ _08495_/B VGND VGND VPWR VPWR _09388_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07445_ _07455_/A _09183_/B VGND VGND VPWR VPWR _07445_/X sky130_fd_sc_hd__and2_1
XFILLER_149_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07376_ _07401_/A VGND VGND VPWR VPWR _09139_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_109_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09115_ _09134_/B _09115_/B VGND VGND VPWR VPWR _09115_/Y sky130_fd_sc_hd__xnor2_1
X_06327_ _14379_/Q _14423_/D VGND VGND VPWR VPWR _06327_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09046_ _09046_/A VGND VGND VPWR VPWR _12758_/D sky130_fd_sc_hd__clkbuf_1
X_06258_ _06258_/A VGND VGND VPWR VPWR _13974_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold440 hold440/A VGND VGND VPWR VPWR hold440/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_135_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06189_ hold520/A _06189_/B VGND VGND VPWR VPWR _06197_/A sky130_fd_sc_hd__xnor2_1
XFILLER_89_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold451 hold451/A VGND VGND VPWR VPWR hold451/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold462 hold462/A VGND VGND VPWR VPWR hold462/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold473 input1/X VGND VGND VPWR VPWR hold473/X sky130_fd_sc_hd__buf_6
XFILLER_116_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold484 hold12/X VGND VGND VPWR VPWR hold484/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold495 hold11/X VGND VGND VPWR VPWR hold495/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09948_ _13700_/Q VGND VGND VPWR VPWR _09957_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_46_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09879_ _13692_/Q _09878_/A _09855_/X VGND VGND VPWR VPWR _09879_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11910_ _14262_/Q _11465_/X _11918_/S VGND VGND VPWR VPWR _11911_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12890_ _12930_/CLK _12890_/D hold1/X VGND VGND VPWR VPWR _12890_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _11841_/A _12149_/A VGND VGND VPWR VPWR _12095_/B sky130_fd_sc_hd__or2b_4
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ _14598_/CLK _14560_/D VGND VGND VPWR VPWR _14560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11772_ _13559_/Q _11772_/B VGND VGND VPWR VPWR _11773_/A sky130_fd_sc_hd__and2_1
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _12896_/Q _10731_/B VGND VGND VPWR VPWR _10724_/A sky130_fd_sc_hd__and2_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _14250_/CLK _13511_/D VGND VGND VPWR VPWR hold351/A sky130_fd_sc_hd__dfxtp_1
X_14491_ _14492_/CLK _14491_/D VGND VGND VPWR VPWR _14491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10654_ _10654_/A VGND VGND VPWR VPWR _12680_/D sky130_fd_sc_hd__clkbuf_1
X_13442_ _13598_/CLK _13442_/D repeater56/X VGND VGND VPWR VPWR _13442_/Q sky130_fd_sc_hd__dfrtp_1
X_13373_ _13377_/CLK _13373_/D repeater57/X VGND VGND VPWR VPWR _13373_/Q sky130_fd_sc_hd__dfrtp_1
X_10585_ _13284_/Q _13035_/Q _13033_/Q _06874_/X VGND VGND VPWR VPWR _13284_/D sky130_fd_sc_hd__o31a_1
XFILLER_154_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12324_ _14577_/Q _12013_/X _12324_/S VGND VGND VPWR VPWR _12325_/A sky130_fd_sc_hd__mux2_1
X_12255_ _11320_/X _14543_/Q _12259_/S VGND VGND VPWR VPWR _12256_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11206_ _13336_/Q _11150_/X _11199_/X _11205_/Y VGND VGND VPWR VPWR _13336_/D sky130_fd_sc_hd__o22a_1
XFILLER_123_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12186_ _14504_/Q _12000_/X _12194_/S VGND VGND VPWR VPWR _12187_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11137_ _11208_/A VGND VGND VPWR VPWR _11137_/X sky130_fd_sc_hd__buf_4
XFILLER_123_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11068_ _14304_/Q _14474_/Q _14230_/Q _14060_/Q _11066_/X _11067_/X VGND VGND VPWR
+ VPWR _11068_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10019_ _10019_/A VGND VGND VPWR VPWR _13910_/D sky130_fd_sc_hd__inv_2
XFILLER_49_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13709_ _14212_/CLK hold351/X VGND VGND VPWR VPWR _13709_/Q sky130_fd_sc_hd__dfxtp_1
X_14689_ _14692_/CLK _14689_/D VGND VGND VPWR VPWR hold191/A sky130_fd_sc_hd__dfxtp_1
X_07230_ _13172_/Q VGND VGND VPWR VPWR _07327_/A sky130_fd_sc_hd__clkbuf_2
X_07161_ _07190_/A _07190_/B VGND VGND VPWR VPWR _07163_/C sky130_fd_sc_hd__and2_1
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06112_ _13941_/D _13942_/D _13943_/D _13964_/D VGND VGND VPWR VPWR _06114_/B sky130_fd_sc_hd__or4_1
XFILLER_8_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07092_ _07093_/A _07093_/B _07093_/C VGND VGND VPWR VPWR _07107_/B sky130_fd_sc_hd__o21a_1
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06043_ hold42/A input20/X _06371_/B _06043_/D VGND VGND VPWR VPWR _06044_/B sky130_fd_sc_hd__and4_1
XFILLER_132_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09802_ _13678_/Q _09802_/B VGND VGND VPWR VPWR _09815_/A sky130_fd_sc_hd__or2_1
X_07994_ _13279_/Q _08001_/B VGND VGND VPWR VPWR _07998_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06945_ _07909_/A VGND VGND VPWR VPWR _06945_/X sky130_fd_sc_hd__buf_2
X_09733_ _14440_/Q _14219_/Q _09836_/B VGND VGND VPWR VPWR _09819_/B sky130_fd_sc_hd__mux2_1
XFILLER_55_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06876_ _06876_/A _06876_/B VGND VGND VPWR VPWR _06877_/B sky130_fd_sc_hd__nor2_1
X_09664_ _14212_/Q _14211_/Q _09731_/A VGND VGND VPWR VPWR _09664_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08615_ _08665_/A _09440_/B _09440_/C VGND VGND VPWR VPWR _08615_/X sky130_fd_sc_hd__and3_1
X_09595_ _09595_/A VGND VGND VPWR VPWR _12812_/D sky130_fd_sc_hd__clkbuf_2
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _08579_/S _13473_/Q VGND VGND VPWR VPWR _08546_/Y sky130_fd_sc_hd__nor2_2
XFILLER_35_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08477_ _13437_/Q _08478_/A VGND VGND VPWR VPWR _08477_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07428_ _07428_/A _07428_/B VGND VGND VPWR VPWR _07428_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07359_ _07396_/A _07364_/A _07359_/C VGND VGND VPWR VPWR _07359_/X sky130_fd_sc_hd__and3_1
XFILLER_164_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10370_ _14211_/D _10374_/A VGND VGND VPWR VPWR _10376_/C sky130_fd_sc_hd__and2_1
XFILLER_164_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09029_ _13215_/Q _13444_/Q _09029_/S VGND VGND VPWR VPWR _09030_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12040_ _12040_/A VGND VGND VPWR VPWR _14409_/D sky130_fd_sc_hd__inv_2
Xhold270 hold270/A VGND VGND VPWR VPWR hold270/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold281 hold281/A VGND VGND VPWR VPWR hold281/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold292 hold292/A VGND VGND VPWR VPWR hold292/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13991_ _14713_/CLK _13991_/D VGND VGND VPWR VPWR _13991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _13274_/CLK _12942_/D VGND VGND VPWR VPWR hold247/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _14179_/CLK _12873_/D VGND VGND VPWR VPWR hold228/A sky130_fd_sc_hd__dfxtp_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _14733_/CLK _14612_/D VGND VGND VPWR VPWR _14612_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _13582_/Q _11828_/B VGND VGND VPWR VPWR _11825_/A sky130_fd_sc_hd__and2_1
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _14543_/CLK _14543_/D VGND VGND VPWR VPWR _14543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _11755_/A VGND VGND VPWR VPWR _14068_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10706_ _10706_/A VGND VGND VPWR VPWR _12931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14474_ _14495_/CLK _14474_/D VGND VGND VPWR VPWR _14474_/Q sky130_fd_sc_hd__dfxtp_1
X_11686_ _11686_/A VGND VGND VPWR VPWR _14025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13425_ _14679_/CLK hold115/X VGND VGND VPWR VPWR _13425_/Q sky130_fd_sc_hd__dfxtp_1
X_10637_ _13814_/Q _14638_/Q VGND VGND VPWR VPWR _13781_/D sky130_fd_sc_hd__xor2_1
XFILLER_10_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10568_ _12991_/D _10566_/X _10575_/A _10558_/B VGND VGND VPWR VPWR _10570_/C sky130_fd_sc_hd__a31oi_1
X_13356_ _13362_/CLK _13356_/D repeater56/X VGND VGND VPWR VPWR _13356_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_6_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12307_ _14569_/Q _11988_/X _12313_/S VGND VGND VPWR VPWR _12308_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13287_ _13525_/CLK hold233/X VGND VGND VPWR VPWR _13287_/Q sky130_fd_sc_hd__dfxtp_1
X_10499_ _10503_/B _10499_/B VGND VGND VPWR VPWR _10500_/A sky130_fd_sc_hd__and2_1
XFILLER_5_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12238_ _12238_/A VGND VGND VPWR VPWR _14535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12169_ _12169_/A VGND VGND VPWR VPWR _14496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 data_i[13] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_4
X_06730_ _06730_/A _06730_/B VGND VGND VPWR VPWR _06731_/B sky130_fd_sc_hd__and2_1
XFILLER_37_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06661_ _06661_/A _06661_/B VGND VGND VPWR VPWR _06661_/X sky130_fd_sc_hd__xor2_1
XFILLER_80_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08400_ _13096_/Q _13377_/Q _08406_/S VGND VGND VPWR VPWR _08401_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09380_ _13592_/Q _09388_/B VGND VGND VPWR VPWR _09382_/A sky130_fd_sc_hd__or2_1
XFILLER_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06592_ _06595_/B _06598_/D VGND VGND VPWR VPWR _06593_/A sky130_fd_sc_hd__and2_1
XFILLER_80_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08331_ _08331_/A _08331_/B VGND VGND VPWR VPWR _08333_/A sky130_fd_sc_hd__and2_1
X_08262_ _10304_/A _08262_/B _08279_/D VGND VGND VPWR VPWR _08268_/B sky130_fd_sc_hd__and3_1
X_14758__69 VGND VGND VPWR VPWR _14758__69/HI _13702_/D sky130_fd_sc_hd__conb_1
X_07213_ _07163_/C _07206_/A _07203_/C _07203_/B VGND VGND VPWR VPWR _07214_/B sky130_fd_sc_hd__o211a_1
X_08193_ _08193_/A _08193_/B VGND VGND VPWR VPWR _08193_/X sky130_fd_sc_hd__xor2_1
XFILLER_118_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07144_ _07144_/A _07144_/B VGND VGND VPWR VPWR _07171_/B sky130_fd_sc_hd__xnor2_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07075_ _07075_/A _07075_/B VGND VGND VPWR VPWR _07077_/C sky130_fd_sc_hd__xor2_1
XFILLER_160_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06026_ _14687_/Q _14683_/Q _14685_/Q VGND VGND VPWR VPWR _06027_/C sky130_fd_sc_hd__or3_1
XFILLER_133_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07977_ _13276_/Q _07981_/B VGND VGND VPWR VPWR _07986_/A sky130_fd_sc_hd__xor2_1
XFILLER_102_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09716_ _09735_/A _09809_/B _09736_/A VGND VGND VPWR VPWR _09720_/B sky130_fd_sc_hd__a21o_1
XFILLER_74_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06928_ _06951_/A _06928_/B VGND VGND VPWR VPWR _06932_/B sky130_fd_sc_hd__nor2_1
XFILLER_142_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09647_ _13419_/Q _13617_/Q _09653_/S VGND VGND VPWR VPWR _09648_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06859_ _06859_/A _07902_/B VGND VGND VPWR VPWR _06859_/X sky130_fd_sc_hd__and2_1
XFILLER_82_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _09579_/B _09579_/C _09579_/A VGND VGND VPWR VPWR _09578_/X sky130_fd_sc_hd__a21o_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08529_ _08529_/A VGND VGND VPWR VPWR _08530_/A sky130_fd_sc_hd__inv_2
XFILLER_70_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11540_ _11540_/A VGND VGND VPWR VPWR _13853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11471_ _11471_/A VGND VGND VPWR VPWR _13825_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10422_ _10426_/B _10422_/B VGND VGND VPWR VPWR _14218_/D sky130_fd_sc_hd__nor2_1
X_13210_ _13593_/CLK hold75/X VGND VGND VPWR VPWR _13210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14190_ _14693_/CLK _14190_/D VGND VGND VPWR VPWR _14190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13141_ _13532_/CLK _13141_/D repeater56/X VGND VGND VPWR VPWR _13141_/Q sky130_fd_sc_hd__dfrtp_1
X_10353_ _13109_/D _13121_/D _10352_/B VGND VGND VPWR VPWR _10353_/X sky130_fd_sc_hd__a21bo_1
XFILLER_125_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13072_ _13294_/CLK _13072_/D VGND VGND VPWR VPWR hold245/A sky130_fd_sc_hd__dfxtp_1
X_10284_ _10284_/A VGND VGND VPWR VPWR _12665_/D sky130_fd_sc_hd__clkbuf_1
X_12023_ _14317_/Q _12022_/X _12026_/S VGND VGND VPWR VPWR _12024_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13974_ _14179_/CLK _13974_/D VGND VGND VPWR VPWR _13974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12925_ _13263_/CLK _12925_/D VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _13686_/CLK _12856_/D VGND VGND VPWR VPWR hold68/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11807_ _11807_/A VGND VGND VPWR VPWR _14096_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _13303_/CLK _12787_/D VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__dfxtp_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _14555_/CLK _14526_/D VGND VGND VPWR VPWR _14526_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11738_ _11749_/A VGND VGND VPWR VPWR _11747_/S sky130_fd_sc_hd__buf_2
XFILLER_119_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14457_ _14733_/CLK _14457_/D VGND VGND VPWR VPWR _14457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11669_ _11691_/A VGND VGND VPWR VPWR _11678_/S sky130_fd_sc_hd__buf_2
X_13408_ _13606_/CLK hold63/X VGND VGND VPWR VPWR _13408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14388_ _14413_/CLK _14388_/D VGND VGND VPWR VPWR _14388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13339_ _14579_/CLK _13339_/D VGND VGND VPWR VPWR _13339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07900_ _06976_/X _07899_/Y _06849_/X VGND VGND VPWR VPWR _13265_/D sky130_fd_sc_hd__a21o_1
XFILLER_102_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08880_ _08881_/A _08881_/B _08881_/C VGND VGND VPWR VPWR _08895_/B sky130_fd_sc_hd__o21a_1
XFILLER_96_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07831_ _07831_/A VGND VGND VPWR VPWR _13256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07762_ _07778_/A _07762_/B VGND VGND VPWR VPWR _07764_/C sky130_fd_sc_hd__nand2_1
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09501_ _09437_/X _09505_/B _09500_/Y _08764_/X VGND VGND VPWR VPWR _13607_/D sky130_fd_sc_hd__a31o_1
XFILLER_65_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06713_ _06712_/A _06712_/C _06712_/B VGND VGND VPWR VPWR _06714_/C sky130_fd_sc_hd__o21ai_1
X_07693_ _07693_/A _07693_/B VGND VGND VPWR VPWR _07695_/A sky130_fd_sc_hd__nor2_1
XFILLER_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09432_ _09447_/A _09447_/C VGND VGND VPWR VPWR _09446_/C sky130_fd_sc_hd__nor2_1
X_06644_ _13353_/Q _13351_/Q _13037_/Q VGND VGND VPWR VPWR _06841_/B sky130_fd_sc_hd__mux2_1
XFILLER_80_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06575_ _12892_/Q _06574_/X _06586_/A VGND VGND VPWR VPWR _06575_/Y sky130_fd_sc_hd__a21oi_1
X_09363_ _13317_/Q _13555_/Q _10822_/A VGND VGND VPWR VPWR _09364_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08314_ _13376_/Q _08314_/B _08317_/D VGND VGND VPWR VPWR _08316_/A sky130_fd_sc_hd__and3_1
X_09294_ _09294_/A VGND VGND VPWR VPWR _12775_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_10 hold42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 input26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 _13340_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08245_ _08245_/A VGND VGND VPWR VPWR _08245_/Y sky130_fd_sc_hd__inv_2
XANTENNA_54 input7/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_65 _13542_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _11115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 hold481/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08176_ _08176_/A VGND VGND VPWR VPWR _08261_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07127_ _07098_/A _07098_/B _07126_/Y VGND VGND VPWR VPWR _07128_/C sky130_fd_sc_hd__o21ai_1
XFILLER_137_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07058_ _07051_/B _07058_/B VGND VGND VPWR VPWR _07077_/A sky130_fd_sc_hd__and2b_1
XFILLER_133_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06009_ _13583_/Q _13584_/Q _13585_/Q _13586_/Q VGND VGND VPWR VPWR _06012_/A sky130_fd_sc_hd__and4_1
XFILLER_102_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10971_ _14598_/Q _14560_/Q _14491_/Q _14443_/Q _10969_/X _10970_/X VGND VGND VPWR
+ VPWR _10972_/A sky130_fd_sc_hd__mux4_1
XFILLER_55_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12710_ _14012_/CLK _12710_/D VGND VGND VPWR VPWR hold431/A sky130_fd_sc_hd__dfxtp_1
X_13690_ _13698_/CLK _13690_/D repeater57/X VGND VGND VPWR VPWR _13690_/Q sky130_fd_sc_hd__dfrtp_1
X_12641_ _12641_/A _12641_/B VGND VGND VPWR VPWR _12642_/A sky130_fd_sc_hd__and2_1
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12572_ _12568_/Y _14739_/Q _12621_/A _12569_/Y _12571_/X VGND VGND VPWR VPWR _12572_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_157_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14311_ _14733_/CLK _14311_/D VGND VGND VPWR VPWR _14311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11523_ _13842_/Q _11522_/X _11523_/S VGND VGND VPWR VPWR _11524_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14242_ _14617_/CLK _14242_/D VGND VGND VPWR VPWR _14242_/Q sky130_fd_sc_hd__dfxtp_1
X_11454_ _13820_/Q _11453_/X _11463_/S VGND VGND VPWR VPWR _11455_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10405_ _10405_/A _10405_/B VGND VGND VPWR VPWR _10405_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_109_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14173_ _14196_/CLK _14173_/D VGND VGND VPWR VPWR _14173_/Q sky130_fd_sc_hd__dfxtp_1
X_11385_ _11444_/B VGND VGND VPWR VPWR _11394_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13124_ _14645_/CLK _13706_/Q VGND VGND VPWR VPWR hold71/A sky130_fd_sc_hd__dfxtp_2
X_10336_ _13109_/Q _13242_/D _10335_/X VGND VGND VPWR VPWR _13167_/D sky130_fd_sc_hd__o21a_1
XFILLER_152_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_9_0_clk clkbuf_4_9_0_clk/A VGND VGND VPWR VPWR clkbuf_4_9_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _10263_/X _10266_/X _10269_/S VGND VGND VPWR VPWR _10268_/A sky130_fd_sc_hd__mux2_1
X_13055_ _13565_/CLK _13055_/D VGND VGND VPWR VPWR hold145/A sky130_fd_sc_hd__dfxtp_1
XFILLER_121_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12006_ _12006_/A VGND VGND VPWR VPWR _14311_/D sky130_fd_sc_hd__clkbuf_1
X_10198_ _14401_/Q _14393_/Q _10627_/A VGND VGND VPWR VPWR _10198_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13957_ _13963_/CLK _13957_/D VGND VGND VPWR VPWR _13957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12908_ _13265_/CLK _12908_/D repeater59/X VGND VGND VPWR VPWR _12908_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13888_ _14050_/CLK _13895_/Q VGND VGND VPWR VPWR _13888_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12839_ _13619_/CLK _12839_/D VGND VGND VPWR VPWR hold61/A sky130_fd_sc_hd__dfxtp_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06360_ _06360_/A VGND VGND VPWR VPWR _14595_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14509_ _14617_/CLK _14509_/D VGND VGND VPWR VPWR _14509_/Q sky130_fd_sc_hd__dfxtp_1
X_06291_ _06291_/A VGND VGND VPWR VPWR _14206_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08030_ hold23/A VGND VGND VPWR VPWR _10803_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_128_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09981_ _09991_/S VGND VGND VPWR VPWR _10596_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_88_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08932_ _08932_/A _08932_/B VGND VGND VPWR VPWR _08959_/B sky130_fd_sc_hd__xnor2_1
XFILLER_115_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08863_ _08863_/A _08863_/B VGND VGND VPWR VPWR _08865_/C sky130_fd_sc_hd__xor2_1
XFILLER_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07814_ _13254_/Q _07821_/B VGND VGND VPWR VPWR _07815_/C sky130_fd_sc_hd__nand2_1
X_08794_ _08789_/A _08790_/X _08793_/Y VGND VGND VPWR VPWR _08794_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_72_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07745_ _07745_/A _07745_/B _07745_/C VGND VGND VPWR VPWR _07746_/B sky130_fd_sc_hd__and3_1
XFILLER_38_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07676_ _07689_/B _07689_/C VGND VGND VPWR VPWR _07677_/B sky130_fd_sc_hd__nor2_1
X_09415_ _09414_/B _09414_/C _13597_/Q VGND VGND VPWR VPWR _09447_/B sky130_fd_sc_hd__a21oi_1
X_06627_ _07214_/A VGND VGND VPWR VPWR _07209_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09346_ _13309_/Q _13547_/Q _09354_/S VGND VGND VPWR VPWR _09347_/A sky130_fd_sc_hd__mux2_1
X_06558_ _06535_/A _06547_/A _06547_/B VGND VGND VPWR VPWR _06558_/X sky130_fd_sc_hd__o21ba_1
XFILLER_40_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09277_ _13552_/Q _09277_/B VGND VGND VPWR VPWR _09277_/X sky130_fd_sc_hd__or2_1
X_06489_ _06488_/Y _06477_/B _06493_/A VGND VGND VPWR VPWR _06490_/B sky130_fd_sc_hd__o21ba_1
XFILLER_138_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08228_ _08126_/X _08270_/B _08228_/S VGND VGND VPWR VPWR _08231_/B sky130_fd_sc_hd__mux2_1
XFILLER_106_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08159_ _08162_/B VGND VGND VPWR VPWR _08177_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11170_ _14311_/Q _14481_/Q _14237_/Q _14067_/Q _11137_/X _11138_/X VGND VGND VPWR
+ VPWR _11170_/X sky130_fd_sc_hd__mux4_1
XFILLER_164_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10121_ _06156_/X _06293_/X _10121_/S VGND VGND VPWR VPWR _10122_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10052_ _10052_/A _13928_/Q VGND VGND VPWR VPWR _10062_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13811_ _13811_/CLK _13811_/D VGND VGND VPWR VPWR _13811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13742_ _13811_/CLK hold434/X VGND VGND VPWR VPWR _13742_/Q sky130_fd_sc_hd__dfxtp_1
X_10954_ _12566_/A VGND VGND VPWR VPWR _12649_/B sky130_fd_sc_hd__buf_2
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13673_ _13673_/CLK _13673_/D repeater56/X VGND VGND VPWR VPWR _13673_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_191_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _14617_/CLK sky130_fd_sc_hd__clkbuf_16
X_10885_ _13159_/Q _10885_/B VGND VGND VPWR VPWR _10886_/A sky130_fd_sc_hd__and2_1
XFILLER_43_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12624_ _14734_/Q _12616_/B _12623_/X _12617_/X VGND VGND VPWR VPWR _14739_/D sky130_fd_sc_hd__o211a_1
XFILLER_157_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12555_ _12555_/A VGND VGND VPWR VPWR _14722_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11506_ _11506_/A VGND VGND VPWR VPWR _13836_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12486_ input28/X VGND VGND VPWR VPWR _12496_/A sky130_fd_sc_hd__clkbuf_2
X_14225_ _14535_/CLK _14225_/D VGND VGND VPWR VPWR _14225_/Q sky130_fd_sc_hd__dfxtp_1
X_11437_ _11437_/A VGND VGND VPWR VPWR _13809_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14156_ _14208_/CLK _14156_/D VGND VGND VPWR VPWR hold67/A sky130_fd_sc_hd__dfxtp_1
X_11368_ _13894_/Q _11362_/X _11364_/B VGND VGND VPWR VPWR _11368_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ _14633_/CLK _13107_/D VGND VGND VPWR VPWR _13107_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _13747_/Q _13107_/Q VGND VGND VPWR VPWR _10321_/C sky130_fd_sc_hd__xnor2_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _14098_/CLK _14087_/D VGND VGND VPWR VPWR _14087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _13760_/Q _11297_/X _11311_/S VGND VGND VPWR VPWR _11300_/A sky130_fd_sc_hd__mux2_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _13039_/CLK _13038_/D VGND VGND VPWR VPWR _13038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07530_ _07530_/A _07530_/B _07530_/C VGND VGND VPWR VPWR _07530_/X sky130_fd_sc_hd__or3_1
XFILLER_34_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07461_ _07461_/A _07461_/B _07461_/C VGND VGND VPWR VPWR _07481_/A sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_182_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _14703_/CLK sky130_fd_sc_hd__clkbuf_16
X_09200_ _13540_/Q _09207_/B VGND VGND VPWR VPWR _09201_/B sky130_fd_sc_hd__or2_1
X_06412_ _14439_/Q _06458_/S VGND VGND VPWR VPWR _06554_/B sky130_fd_sc_hd__and2_1
X_07392_ _13139_/Q _09130_/B _07381_/A VGND VGND VPWR VPWR _07415_/B sky130_fd_sc_hd__a21oi_1
XFILLER_31_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06343_ _14108_/Q _14092_/Q _06345_/S VGND VGND VPWR VPWR _06344_/A sky130_fd_sc_hd__mux2_1
X_09131_ _13530_/Q _09126_/B _07356_/B _13529_/Q VGND VGND VPWR VPWR _09131_/X sky130_fd_sc_hd__o211a_1
XFILLER_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09062_ _13229_/Q _13458_/Q _09064_/S VGND VGND VPWR VPWR _09063_/A sky130_fd_sc_hd__mux2_1
X_06274_ _06274_/A VGND VGND VPWR VPWR _13955_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08013_ _08013_/A _08013_/B _08007_/Y _08008_/X VGND VGND VPWR VPWR _08018_/C sky130_fd_sc_hd__or4bb_1
XFILLER_163_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09964_ _13505_/Q _13694_/Q _09968_/S VGND VGND VPWR VPWR _09965_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08915_ _08886_/A _08886_/B _08914_/Y VGND VGND VPWR VPWR _08916_/C sky130_fd_sc_hd__o21ai_1
XFILLER_98_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ _09895_/A VGND VGND VPWR VPWR _13696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08846_ _08839_/B _08846_/B VGND VGND VPWR VPWR _08865_/A sky130_fd_sc_hd__and2b_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08777_ _08786_/A _08786_/B _08542_/A VGND VGND VPWR VPWR _08777_/X sky130_fd_sc_hd__a21o_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05989_ _14107_/Q _14108_/Q _14109_/Q VGND VGND VPWR VPWR _05992_/A sky130_fd_sc_hd__and3_1
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ _07753_/B _07728_/B VGND VGND VPWR VPWR _07729_/B sky130_fd_sc_hd__xnor2_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07659_ _07659_/A _07659_/B _07659_/C VGND VGND VPWR VPWR _07660_/B sky130_fd_sc_hd__or3_1
XFILLER_26_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_173_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _14737_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10670_ _14341_/Q _10671_/C _10669_/Y VGND VGND VPWR VPWR _12916_/D sky130_fd_sc_hd__a21oi_1
XFILLER_138_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09329_ _09329_/A VGND VGND VPWR VPWR _12791_/D sky130_fd_sc_hd__clkbuf_1
X_12340_ _14642_/Q _12340_/B VGND VGND VPWR VPWR _12341_/A sky130_fd_sc_hd__and2_1
XFILLER_138_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12271_ _12271_/A VGND VGND VPWR VPWR _14550_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14010_ _14010_/CLK _14010_/D VGND VGND VPWR VPWR _14010_/Q sky130_fd_sc_hd__dfxtp_1
X_11222_ _14033_/Q _13999_/Q _13839_/Q _14551_/Q _10993_/A _10995_/A VGND VGND VPWR
+ VPWR _11223_/A sky130_fd_sc_hd__mux4_1
XFILLER_135_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11153_ _11153_/A VGND VGND VPWR VPWR _11153_/X sky130_fd_sc_hd__buf_2
XFILLER_122_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10104_ _10139_/A _14145_/Q VGND VGND VPWR VPWR _10143_/A sky130_fd_sc_hd__xnor2_1
X_11084_ _11155_/A VGND VGND VPWR VPWR _11084_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10035_ _10035_/A VGND VGND VPWR VPWR _13971_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11986_ _14305_/Q _11984_/X _11998_/S VGND VGND VPWR VPWR _11987_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13725_ _13727_/CLK hold279/X VGND VGND VPWR VPWR _13725_/Q sky130_fd_sc_hd__dfxtp_1
X_10937_ _14596_/Q _14558_/Q _14489_/Q _14441_/Q _11208_/A _11209_/A VGND VGND VPWR
+ VPWR _10938_/A sky130_fd_sc_hd__mux4_1
XFILLER_17_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_164_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _14555_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13656_ _13657_/CLK _13656_/D VGND VGND VPWR VPWR _13656_/Q sky130_fd_sc_hd__dfxtp_1
X_10868_ _13151_/Q _10874_/B VGND VGND VPWR VPWR _10869_/A sky130_fd_sc_hd__and2_1
XFILLER_13_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12607_ _12607_/A VGND VGND VPWR VPWR _14732_/D sky130_fd_sc_hd__clkbuf_1
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13587_ _13587_/CLK hold222/X VGND VGND VPWR VPWR hold173/A sky130_fd_sc_hd__dfxtp_2
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10799_ _13020_/Q _10801_/B VGND VGND VPWR VPWR _10800_/A sky130_fd_sc_hd__and2_1
X_12538_ _12538_/A VGND VGND VPWR VPWR _14714_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12469_ _12469_/A VGND VGND VPWR VPWR _14665_/D sky130_fd_sc_hd__clkbuf_1
X_14208_ _14208_/CLK _14208_/D VGND VGND VPWR VPWR _14208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14139_ _14716_/CLK _14139_/D VGND VGND VPWR VPWR hold330/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06961_ _08002_/B VGND VGND VPWR VPWR _08015_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_39_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08700_ _09524_/B VGND VGND VPWR VPWR _09511_/B sky130_fd_sc_hd__clkbuf_2
X_05912_ _06091_/A VGND VGND VPWR VPWR _06273_/S sky130_fd_sc_hd__clkinv_2
X_09680_ _09758_/A _09679_/C _13668_/Q VGND VGND VPWR VPWR _09680_/X sky130_fd_sc_hd__a21o_1
X_06892_ _07989_/B VGND VGND VPWR VPWR _08001_/B sky130_fd_sc_hd__clkbuf_2
X_08631_ _08665_/A _09450_/B VGND VGND VPWR VPWR _08631_/X sky130_fd_sc_hd__and2_1
XFILLER_94_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08562_ _08556_/B _08561_/Y _09404_/S VGND VGND VPWR VPWR _08563_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07513_ _13152_/Q _07513_/B VGND VGND VPWR VPWR _07515_/A sky130_fd_sc_hd__nand2_1
XFILLER_120_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_155_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _14712_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08493_ _08567_/A _08497_/B VGND VGND VPWR VPWR _08495_/B sky130_fd_sc_hd__and2b_1
X_07444_ _07444_/A VGND VGND VPWR VPWR _09183_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07375_ _07375_/A _07375_/B _07375_/C VGND VGND VPWR VPWR _07401_/A sky130_fd_sc_hd__nand3_2
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09114_ _09114_/A _09134_/A VGND VGND VPWR VPWR _09115_/B sky130_fd_sc_hd__nand2_1
X_06326_ _06324_/A _06324_/Y _14414_/D _06325_/X VGND VGND VPWR VPWR _14424_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06257_ _06256_/X _06076_/A _06257_/S VGND VGND VPWR VPWR _06258_/A sky130_fd_sc_hd__mux2_1
X_09045_ _13222_/Q _13451_/Q _09051_/S VGND VGND VPWR VPWR _09046_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06188_ _14424_/Q _14422_/Q _14426_/Q VGND VGND VPWR VPWR _06189_/B sky130_fd_sc_hd__mux2_1
Xhold430 hold430/A VGND VGND VPWR VPWR hold430/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold441 hold441/A VGND VGND VPWR VPWR hold441/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold452 hold452/A VGND VGND VPWR VPWR hold452/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold463 hold463/A VGND VGND VPWR VPWR hold463/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold474 hold474/A VGND VGND VPWR VPWR hold474/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold485 hold485/A VGND VGND VPWR VPWR hold485/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_145_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold496 hold496/A VGND VGND VPWR VPWR hold496/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_131_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09947_ _09947_/A VGND VGND VPWR VPWR _12860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _09878_/A _09878_/B VGND VGND VPWR VPWR _13691_/D sky130_fd_sc_hd__nor2_1
XFILLER_38_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08829_ _13430_/Q VGND VGND VPWR VPWR _08929_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _11840_/A VGND VGND VPWR VPWR _14192_/D sky130_fd_sc_hd__inv_2
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_146_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _14608_/CLK sky130_fd_sc_hd__clkbuf_16
X_11771_ _11771_/A VGND VGND VPWR VPWR _14080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _13704_/CLK hold268/X VGND VGND VPWR VPWR _13510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10722_ _13031_/D VGND VGND VPWR VPWR _10731_/B sky130_fd_sc_hd__clkbuf_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _14619_/CLK _14490_/D VGND VGND VPWR VPWR _14490_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13441_ _13702_/CLK _13441_/D repeater56/X VGND VGND VPWR VPWR _13441_/Q sky130_fd_sc_hd__dfrtp_1
X_10653_ _13713_/Q _11382_/B VGND VGND VPWR VPWR _10654_/A sky130_fd_sc_hd__and2_1
XFILLER_155_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13372_ _13372_/CLK _13372_/D repeater57/X VGND VGND VPWR VPWR _13372_/Q sky130_fd_sc_hd__dfrtp_1
X_10584_ _13168_/Q hold487/X _13163_/Q _07343_/X VGND VGND VPWR VPWR _13163_/D sky130_fd_sc_hd__o31a_1
XFILLER_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12323_ _12323_/A VGND VGND VPWR VPWR _14576_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12254_ _12254_/A VGND VGND VPWR VPWR _14542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11205_ _11242_/A _11205_/B VGND VGND VPWR VPWR _11205_/Y sky130_fd_sc_hd__nand2_1
X_12185_ _12185_/A VGND VGND VPWR VPWR _12194_/S sky130_fd_sc_hd__buf_2
X_11136_ _11207_/A VGND VGND VPWR VPWR _11136_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11067_ _11209_/A VGND VGND VPWR VPWR _11067_/X sky130_fd_sc_hd__buf_2
XFILLER_76_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10018_ _10056_/A VGND VGND VPWR VPWR _14038_/D sky130_fd_sc_hd__inv_2
XFILLER_76_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11969_ _12001_/A VGND VGND VPWR VPWR _11982_/S sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_137_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _14294_/CLK sky130_fd_sc_hd__clkbuf_16
X_13708_ _14645_/CLK _13708_/D VGND VGND VPWR VPWR _13708_/Q sky130_fd_sc_hd__dfxtp_1
X_14688_ _14688_/CLK hold96/X VGND VGND VPWR VPWR _14688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13639_ _14327_/CLK hold407/X VGND VGND VPWR VPWR _13639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07160_ _07163_/B VGND VGND VPWR VPWR _07203_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_9_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06111_ _06109_/X _06110_/X _11593_/B VGND VGND VPWR VPWR _13964_/D sky130_fd_sc_hd__o21a_1
XFILLER_9_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07091_ _14634_/Q _13115_/D VGND VGND VPWR VPWR _07093_/C sky130_fd_sc_hd__nand2_1
XFILLER_133_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06042_ input17/X input21/X input22/X VGND VGND VPWR VPWR _06043_/D sky130_fd_sc_hd__and3_1
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09801_ _13678_/Q _09802_/B VGND VGND VPWR VPWR _09803_/A sky130_fd_sc_hd__and2_1
XFILLER_115_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07993_ _06793_/A _07995_/B _07992_/Y _07940_/X VGND VGND VPWR VPWR _13278_/D sky130_fd_sc_hd__a31o_1
XFILLER_140_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09732_ _14217_/Q _14215_/Q _09836_/B VGND VGND VPWR VPWR _09732_/X sky130_fd_sc_hd__mux2_1
X_06944_ _06861_/X _06942_/Y _06943_/X _06907_/X VGND VGND VPWR VPWR _13020_/D sky130_fd_sc_hd__a31o_1
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09663_ _13709_/Q VGND VGND VPWR VPWR _09731_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06875_ _13011_/Q _07895_/B _07895_/C VGND VGND VPWR VPWR _06877_/A sky130_fd_sc_hd__nand3_1
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08614_ _08614_/A _08614_/B VGND VGND VPWR VPWR _08614_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_54_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09594_ _13395_/Q _13593_/Q _09598_/S VGND VGND VPWR VPWR _09595_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08545_ _13473_/Q _14256_/Q _08545_/S VGND VGND VPWR VPWR _08545_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_128_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _13972_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08476_ _08490_/A _08490_/B VGND VGND VPWR VPWR _08478_/A sky130_fd_sc_hd__xor2_1
XFILLER_23_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07427_ _07411_/X _07424_/X _07425_/Y _07426_/X VGND VGND VPWR VPWR _13143_/D sky130_fd_sc_hd__a31o_1
X_07358_ _07358_/A _07358_/B VGND VGND VPWR VPWR _07358_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_109_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06309_ _13875_/Q _13859_/Q _06309_/S VGND VGND VPWR VPWR _06310_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07289_ _13134_/Q _09098_/B VGND VGND VPWR VPWR _07305_/A sky130_fd_sc_hd__nor2_1
X_09028_ _09028_/A VGND VGND VPWR VPWR _12750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold260 hold260/A VGND VGND VPWR VPWR hold260/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold271 hold271/A VGND VGND VPWR VPWR hold271/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold282 hold282/A VGND VGND VPWR VPWR hold282/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold293 hold293/A VGND VGND VPWR VPWR hold293/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13990_ _14713_/CLK _13990_/D VGND VGND VPWR VPWR _13990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12941_ _12974_/CLK _12941_/D VGND VGND VPWR VPWR hold302/A sky130_fd_sc_hd__dfxtp_1
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12872_ _13698_/CLK _12872_/D VGND VGND VPWR VPWR hold181/A sky130_fd_sc_hd__dfxtp_1
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _14619_/CLK _14611_/D VGND VGND VPWR VPWR _14611_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11823_ _11823_/A VGND VGND VPWR VPWR _14103_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _14075_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _14543_/CLK _14542_/D VGND VGND VPWR VPWR _14542_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _11343_/X _14068_/Q _11758_/S VGND VGND VPWR VPWR _11755_/A sky130_fd_sc_hd__mux2_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _12888_/Q _10709_/B VGND VGND VPWR VPWR _10706_/A sky130_fd_sc_hd__and2_1
XFILLER_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14473_ _14600_/CLK _14473_/D VGND VGND VPWR VPWR _14473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11685_ _14025_/Q _11488_/X _11689_/S VGND VGND VPWR VPWR _11686_/A sky130_fd_sc_hd__mux2_1
X_13424_ _14679_/CLK hold394/X VGND VGND VPWR VPWR _13424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10636_ _10636_/A _13814_/Q VGND VGND VPWR VPWR _13780_/D sky130_fd_sc_hd__xor2_1
XFILLER_127_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13355_ _13657_/CLK _13355_/D hold1/X VGND VGND VPWR VPWR _13355_/Q sky130_fd_sc_hd__dfrtp_1
X_10567_ _10567_/A _10573_/C VGND VGND VPWR VPWR _10575_/A sky130_fd_sc_hd__nand2_1
XFILLER_10_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12306_ _12306_/A VGND VGND VPWR VPWR _14568_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13286_ _13525_/CLK hold119/X VGND VGND VPWR VPWR _13286_/Q sky130_fd_sc_hd__dfxtp_1
X_10498_ _10498_/A _10498_/B _10498_/C VGND VGND VPWR VPWR _10499_/B sky130_fd_sc_hd__nand3_1
X_12237_ _11294_/X _14535_/Q _12237_/S VGND VGND VPWR VPWR _12238_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12168_ _14496_/Q _11975_/X _12172_/S VGND VGND VPWR VPWR _12169_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11119_ _11190_/A VGND VGND VPWR VPWR _11177_/A sky130_fd_sc_hd__clkbuf_4
X_12099_ _12099_/A VGND VGND VPWR VPWR _14465_/D sky130_fd_sc_hd__clkbuf_1
Xinput6 data_i[14] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__buf_6
XFILLER_110_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06660_ _12998_/Q _07807_/B VGND VGND VPWR VPWR _06661_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06591_ _12896_/Q _12897_/Q VGND VGND VPWR VPWR _06598_/D sky130_fd_sc_hd__and2_1
XFILLER_33_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08330_ _13381_/Q VGND VGND VPWR VPWR _08331_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_32_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08261_ _08261_/A VGND VGND VPWR VPWR _10304_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07212_ _07207_/A _07206_/B _07208_/B _07208_/A VGND VGND VPWR VPWR _07215_/A sky130_fd_sc_hd__a22o_1
XFILLER_119_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08192_ _08169_/A _08170_/A _08169_/B _08180_/Y _08191_/Y VGND VGND VPWR VPWR _08193_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_119_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07143_ _07165_/A _07190_/B VGND VGND VPWR VPWR _07144_/B sky130_fd_sc_hd__nand2_1
XFILLER_146_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07074_ _07074_/A _07074_/B VGND VGND VPWR VPWR _07075_/B sky130_fd_sc_hd__or2_1
XFILLER_145_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06025_ _14686_/Q _06025_/B VGND VGND VPWR VPWR _06353_/A sky130_fd_sc_hd__nand2_1
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07976_ _07925_/A _07973_/X _07975_/Y VGND VGND VPWR VPWR _07987_/A sky130_fd_sc_hd__o21ai_4
XFILLER_142_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09715_ _14220_/Q _14218_/Q _09715_/S VGND VGND VPWR VPWR _09809_/B sky130_fd_sc_hd__mux2_1
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06927_ _06899_/Y _06951_/B _06926_/X VGND VGND VPWR VPWR _06928_/B sky130_fd_sc_hd__o21ba_1
XFILLER_27_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09646_ _09646_/A VGND VGND VPWR VPWR _12835_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06858_ _06858_/A _06876_/A VGND VGND VPWR VPWR _06870_/B sky130_fd_sc_hd__or2_1
XFILLER_27_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _09577_/A _09577_/B VGND VGND VPWR VPWR _09579_/A sky130_fd_sc_hd__nand2_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06789_ _13007_/Q _07863_/B _07863_/C VGND VGND VPWR VPWR _06791_/A sky130_fd_sc_hd__and3_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08528_ _13439_/Q _09394_/B VGND VGND VPWR VPWR _08529_/A sky130_fd_sc_hd__and2_1
X_08459_ _08459_/A _08459_/B VGND VGND VPWR VPWR _08459_/X sky130_fd_sc_hd__xor2_1
X_11470_ _13825_/Q _11469_/X _11479_/S VGND VGND VPWR VPWR _11471_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10421_ _10421_/A _10421_/B _10421_/C VGND VGND VPWR VPWR _10422_/B sky130_fd_sc_hd__nor3_1
XFILLER_136_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13140_ _13532_/CLK _13140_/D hold1/X VGND VGND VPWR VPWR _13140_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10352_ _10352_/A _10352_/B VGND VGND VPWR VPWR _13039_/D sky130_fd_sc_hd__xnor2_1
XFILLER_164_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13071_ _14555_/CLK _13071_/D VGND VGND VPWR VPWR hold162/A sky130_fd_sc_hd__dfxtp_1
X_10283_ _10282_/X _10279_/X _10592_/B VGND VGND VPWR VPWR _10284_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12022_ _12022_/A VGND VGND VPWR VPWR _12022_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13973_ _14179_/CLK _13973_/D VGND VGND VPWR VPWR _13973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12924_ _13263_/CLK _12924_/D VGND VGND VPWR VPWR hold275/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12855_ _13727_/CLK _12855_/D VGND VGND VPWR VPWR hold313/A sky130_fd_sc_hd__dfxtp_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _13574_/Q _11806_/B VGND VGND VPWR VPWR _11807_/A sky130_fd_sc_hd__and2_1
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _13574_/CLK _12786_/D VGND VGND VPWR VPWR hold386/A sky130_fd_sc_hd__dfxtp_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14525_ _14557_/CLK _14525_/D VGND VGND VPWR VPWR _14525_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _11737_/A VGND VGND VPWR VPWR _14060_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14456_ _14619_/CLK _14456_/D VGND VGND VPWR VPWR _14456_/Q sky130_fd_sc_hd__dfxtp_1
X_11668_ _11668_/A VGND VGND VPWR VPWR _14017_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13407_ _13606_/CLK hold444/X VGND VGND VPWR VPWR _13407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10619_ _10119_/S _10616_/X _10617_/X _10618_/X _14166_/Q VGND VGND VPWR VPWR _14208_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14387_ _14413_/CLK _14387_/D VGND VGND VPWR VPWR _14387_/Q sky130_fd_sc_hd__dfxtp_1
X_11599_ _11712_/B VGND VGND VPWR VPWR _12614_/A sky130_fd_sc_hd__inv_2
XFILLER_128_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13338_ _14579_/CLK _13338_/D VGND VGND VPWR VPWR _13338_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_116_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13269_ _13273_/CLK _13269_/D repeater59/X VGND VGND VPWR VPWR _13269_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07830_ _07832_/B _07829_/Y _07843_/S VGND VGND VPWR VPWR _07831_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07761_ _07761_/A _07759_/C VGND VGND VPWR VPWR _07762_/B sky130_fd_sc_hd__or2b_1
XFILLER_2_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09500_ _09500_/A _09500_/B _09509_/C VGND VGND VPWR VPWR _09500_/Y sky130_fd_sc_hd__nand3_1
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06712_ _06712_/A _06712_/B _06712_/C VGND VGND VPWR VPWR _06730_/B sky130_fd_sc_hd__or3_1
X_07692_ _13111_/Q _13112_/Q _07723_/C _14584_/Q VGND VGND VPWR VPWR _07693_/B sky130_fd_sc_hd__and4_1
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09431_ _13599_/Q _09438_/B VGND VGND VPWR VPWR _09454_/B sky130_fd_sc_hd__xnor2_1
XFILLER_64_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06643_ _06643_/A VGND VGND VPWR VPWR _06736_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09362_ _09362_/A VGND VGND VPWR VPWR _12806_/D sky130_fd_sc_hd__clkbuf_1
X_06574_ _06584_/C VGND VGND VPWR VPWR _06574_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_08313_ _13375_/Q _08309_/A _08312_/Y _07239_/X VGND VGND VPWR VPWR _13375_/D sky130_fd_sc_hd__o211a_1
X_09293_ _13285_/Q _13523_/Q _09299_/S VGND VGND VPWR VPWR _09294_/A sky130_fd_sc_hd__mux2_1
XANTENNA_11 hold42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 input26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08244_ _08244_/A _08256_/A VGND VGND VPWR VPWR _08247_/A sky130_fd_sc_hd__or2b_1
XANTENNA_44 _13322_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 input8/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_66 _13547_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_77 _11116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_88 _13700_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08175_ _08176_/A _08262_/B _08177_/A VGND VGND VPWR VPWR _08175_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07126_ _07126_/A _07126_/B VGND VGND VPWR VPWR _07126_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07057_ _07057_/A VGND VGND VPWR VPWR _13344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06008_ hold173/A _13556_/Q _13557_/Q _13558_/Q VGND VGND VPWR VPWR _06008_/X sky130_fd_sc_hd__and4_1
XFILLER_0_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07959_ _07948_/A _07952_/X _07972_/B _06743_/A VGND VGND VPWR VPWR _07959_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_101_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10970_ _11153_/A VGND VGND VPWR VPWR _10970_/X sky130_fd_sc_hd__buf_2
XFILLER_44_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09629_ _13411_/Q _13609_/Q _09631_/S VGND VGND VPWR VPWR _09630_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12640_ _10914_/X _12625_/B _12631_/C VGND VGND VPWR VPWR _12641_/B sky130_fd_sc_hd__a21o_1
XFILLER_71_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12571_ _12569_/Y _12621_/A _12619_/A _12570_/Y VGND VGND VPWR VPWR _12571_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_50_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _13353_/CLK sky130_fd_sc_hd__clkbuf_16
X_14310_ _14667_/CLK _14310_/D VGND VGND VPWR VPWR _14310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11522_ _12025_/A VGND VGND VPWR VPWR _11522_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14241_ _14617_/CLK _14241_/D VGND VGND VPWR VPWR _14241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11453_ _14695_/Q VGND VGND VPWR VPWR _11453_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10404_ _10378_/A _10431_/A _10403_/X VGND VGND VPWR VPWR _10405_/B sky130_fd_sc_hd__o21a_1
X_14172_ _14201_/CLK _14172_/D VGND VGND VPWR VPWR _14172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11384_ _11429_/A VGND VGND VPWR VPWR _11444_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_164_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13123_ _14645_/CLK hold425/X VGND VGND VPWR VPWR hold186/A sky130_fd_sc_hd__dfxtp_2
XFILLER_152_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10335_ _13109_/Q _13242_/D _10334_/B VGND VGND VPWR VPWR _10335_/X sky130_fd_sc_hd__a21bo_1
XFILLER_3_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _13565_/CLK _13054_/D VGND VGND VPWR VPWR hold124/A sky130_fd_sc_hd__dfxtp_1
X_10266_ _10259_/X _14357_/D _10266_/S VGND VGND VPWR VPWR _10266_/X sky130_fd_sc_hd__mux2_1
X_12005_ _14311_/Q _12004_/X _12014_/S VGND VGND VPWR VPWR _12006_/A sky130_fd_sc_hd__mux2_1
X_10197_ _10197_/A VGND VGND VPWR VPWR _10627_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_93_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13956_ _13963_/CLK _13956_/D VGND VGND VPWR VPWR _13956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12907_ _13274_/CLK _12907_/D repeater59/X VGND VGND VPWR VPWR _12907_/Q sky130_fd_sc_hd__dfrtp_1
X_13887_ _14210_/CLK _13887_/D VGND VGND VPWR VPWR hold316/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12838_ _14327_/CLK _12838_/D VGND VGND VPWR VPWR hold401/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _13855_/CLK _12769_/D VGND VGND VPWR VPWR hold274/A sky130_fd_sc_hd__dfxtp_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _13039_/CLK sky130_fd_sc_hd__clkbuf_16
X_06290_ _06289_/X _06146_/A _06290_/S VGND VGND VPWR VPWR _06291_/A sky130_fd_sc_hd__mux2_1
X_14508_ _14579_/CLK _14508_/D VGND VGND VPWR VPWR _14508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput20 input20/A VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__clkbuf_2
X_14439_ _14439_/CLK _14439_/D VGND VGND VPWR VPWR _14439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09980_ _14632_/Q _09980_/B VGND VGND VPWR VPWR _09991_/S sky130_fd_sc_hd__xnor2_1
XFILLER_143_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08931_ _08953_/A _08978_/B VGND VGND VPWR VPWR _08932_/B sky130_fd_sc_hd__nand2_1
XFILLER_130_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08862_ _08862_/A _08862_/B VGND VGND VPWR VPWR _08863_/B sky130_fd_sc_hd__or2_1
X_07813_ _13254_/Q _07813_/B VGND VGND VPWR VPWR _07815_/B sky130_fd_sc_hd__or2_1
XFILLER_96_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08793_ _13466_/Q _09581_/B VGND VGND VPWR VPWR _08793_/Y sky130_fd_sc_hd__xnor2_1
X_07744_ _07745_/A _07785_/C _07745_/C VGND VGND VPWR VPWR _07746_/A sky130_fd_sc_hd__a21oi_1
XFILLER_53_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07675_ _07675_/A _07675_/B _07675_/C VGND VGND VPWR VPWR _07689_/C sky130_fd_sc_hd__nor3_1
XFILLER_26_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09414_ _13597_/Q _09414_/B _09414_/C VGND VGND VPWR VPWR _09447_/A sky130_fd_sc_hd__and3_1
X_06626_ _14631_/Q _13116_/D VGND VGND VPWR VPWR _07214_/A sky130_fd_sc_hd__xor2_4
XFILLER_25_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09345_ _10831_/A VGND VGND VPWR VPWR _09354_/S sky130_fd_sc_hd__clkbuf_2
X_06557_ _06557_/A _06557_/B VGND VGND VPWR VPWR _06567_/A sky130_fd_sc_hd__or2_1
XFILLER_40_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _13304_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09276_ _13552_/Q _09277_/B VGND VGND VPWR VPWR _09276_/Y sky130_fd_sc_hd__nand2_1
X_06488_ _06488_/A VGND VGND VPWR VPWR _06488_/Y sky130_fd_sc_hd__inv_2
X_08227_ _08218_/X _08225_/Y _08226_/Y VGND VGND VPWR VPWR _13363_/D sky130_fd_sc_hd__a21oi_1
XFILLER_5_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08158_ _14012_/Q _14010_/Q _08161_/S VGND VGND VPWR VPWR _08250_/B sky130_fd_sc_hd__mux2_1
X_07109_ _13112_/D _07141_/C _07163_/B hold515/A VGND VGND VPWR VPWR _07111_/A sky130_fd_sc_hd__a22oi_1
XFILLER_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08089_ _12980_/Q _13280_/Q _08095_/S VGND VGND VPWR VPWR _08090_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10120_ _10120_/A VGND VGND VPWR VPWR _14202_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_99_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _13799_/CLK sky130_fd_sc_hd__clkbuf_16
X_10051_ _10051_/A VGND VGND VPWR VPWR _13951_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13810_ _13811_/CLK _13810_/D VGND VGND VPWR VPWR _13810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13741_ _13811_/CLK hold323/X VGND VGND VPWR VPWR _13741_/Q sky130_fd_sc_hd__dfxtp_1
X_10953_ _12645_/A _10950_/X _10952_/X _10929_/X VGND VGND VPWR VPWR _10953_/X sky130_fd_sc_hd__o211a_1
XFILLER_44_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13672_ _13673_/CLK _13672_/D repeater56/X VGND VGND VPWR VPWR _13672_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_44_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10884_ _10884_/A VGND VGND VPWR VPWR _13200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12623_ _14739_/Q _12623_/B VGND VGND VPWR VPWR _12623_/X sky130_fd_sc_hd__or2_1
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _13558_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_156_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12554_ _11354_/X _14722_/Q _12554_/S VGND VGND VPWR VPWR _12555_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11505_ _13836_/Q _11504_/X _11511_/S VGND VGND VPWR VPWR _11506_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12485_ _12485_/A VGND VGND VPWR VPWR _14673_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14224_ _14535_/CLK _14224_/D VGND VGND VPWR VPWR _14224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11436_ _13740_/Q _11438_/B VGND VGND VPWR VPWR _11437_/A sky130_fd_sc_hd__and2_1
XFILLER_138_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14155_ _14294_/CLK hold67/X VGND VGND VPWR VPWR hold383/A sky130_fd_sc_hd__dfxtp_1
X_11367_ _11367_/A VGND VGND VPWR VPWR _13776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13106_ _14633_/CLK _13106_/D VGND VGND VPWR VPWR _13106_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ _10315_/A _10317_/B _10315_/B VGND VGND VPWR VPWR _13471_/D sky130_fd_sc_hd__a21bo_1
X_14086_ _14397_/CLK _14086_/D VGND VGND VPWR VPWR _14086_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _11330_/A VGND VGND VPWR VPWR _11311_/S sky130_fd_sc_hd__buf_2
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _13353_/CLK _13037_/D VGND VGND VPWR VPWR _13037_/Q sky130_fd_sc_hd__dfxtp_1
X_10249_ _14529_/D _10248_/X _14555_/D VGND VGND VPWR VPWR _10250_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13939_ _13978_/CLK _13939_/D VGND VGND VPWR VPWR _13939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07460_ _07424_/X _07434_/A _07442_/B _07454_/C _07459_/X VGND VGND VPWR VPWR _07477_/B
+ sky130_fd_sc_hd__o41ai_4
XFILLER_22_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06411_ _13106_/D VGND VGND VPWR VPWR _06458_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_34_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07391_ _13141_/Q _07395_/A VGND VGND VPWR VPWR _07414_/A sky130_fd_sc_hd__xnor2_1
XFILLER_15_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _14108_/CLK sky130_fd_sc_hd__clkbuf_16
X_09130_ _13531_/Q _09130_/B VGND VGND VPWR VPWR _09161_/A sky130_fd_sc_hd__xnor2_1
X_06342_ _06342_/A VGND VGND VPWR VPWR _14406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09061_ _09061_/A VGND VGND VPWR VPWR _12764_/D sky130_fd_sc_hd__clkbuf_1
X_06273_ _13809_/Q _13793_/Q _06273_/S VGND VGND VPWR VPWR _06274_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08012_ _13280_/Q _13281_/Q _06895_/B VGND VGND VPWR VPWR _08018_/B sky130_fd_sc_hd__o21ai_1
X_09963_ _09963_/A VGND VGND VPWR VPWR _12867_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08914_ _08914_/A _08914_/B VGND VGND VPWR VPWR _08914_/Y sky130_fd_sc_hd__nand2_1
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _09894_/A _09894_/B _09894_/C VGND VGND VPWR VPWR _09895_/A sky130_fd_sc_hd__and3_1
XFILLER_100_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08845_ _08845_/A VGND VGND VPWR VPWR _14247_/D sky130_fd_sc_hd__clkbuf_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08776_ _08786_/A _08786_/B VGND VGND VPWR VPWR _08776_/Y sky130_fd_sc_hd__nor2_1
XFILLER_150_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05988_ hold77/A _14094_/Q _14095_/Q _14098_/Q VGND VGND VPWR VPWR _05993_/C sky130_fd_sc_hd__and4_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07727_ _07693_/A _07695_/B _07693_/B VGND VGND VPWR VPWR _07728_/B sky130_fd_sc_hd__o21ba_1
XFILLER_150_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07658_ _07659_/A _07659_/B _07659_/C VGND VGND VPWR VPWR _07683_/A sky130_fd_sc_hd__o21ai_2
XFILLER_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06609_ _06620_/B _06609_/B _06609_/C VGND VGND VPWR VPWR _06610_/A sky130_fd_sc_hd__and3b_1
XFILLER_80_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_8_0_clk clkbuf_4_9_0_clk/A VGND VGND VPWR VPWR clkbuf_4_8_0_clk/X sky130_fd_sc_hd__clkbuf_2
X_07589_ _07581_/A _07587_/Y _07585_/Y _07586_/X VGND VGND VPWR VPWR _07589_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_9_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09328_ _13301_/Q _13539_/Q _09332_/S VGND VGND VPWR VPWR _09329_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09259_ _09264_/A _09259_/B VGND VGND VPWR VPWR _09267_/A sky130_fd_sc_hd__nand2_1
XFILLER_138_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12270_ _11354_/X _14550_/Q _12270_/S VGND VGND VPWR VPWR _12271_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11221_ _14315_/Q _14485_/Q _14241_/Q _14071_/Q _11208_/X _11209_/X VGND VGND VPWR
+ VPWR _11221_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11152_ _12585_/A VGND VGND VPWR VPWR _11152_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_150_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10103_ _10103_/A VGND VGND VPWR VPWR _14294_/D sky130_fd_sc_hd__inv_2
XFILLER_1_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11083_ _14023_/Q _13989_/Q _13829_/Q _14541_/Q _11081_/X _11082_/X VGND VGND VPWR
+ VPWR _11085_/A sky130_fd_sc_hd__mux4_1
XFILLER_150_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10034_ _06086_/X _06260_/X _10034_/S VGND VGND VPWR VPWR _10035_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11985_ _12001_/A VGND VGND VPWR VPWR _11998_/S sky130_fd_sc_hd__buf_2
XFILLER_16_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10936_ _11153_/A VGND VGND VPWR VPWR _11209_/A sky130_fd_sc_hd__buf_2
X_13724_ _13727_/CLK hold452/X VGND VGND VPWR VPWR _13724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10867_ _10867_/A VGND VGND VPWR VPWR _13192_/D sky130_fd_sc_hd__clkbuf_1
X_13655_ _13657_/CLK _13655_/D VGND VGND VPWR VPWR _13655_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12606_ _12608_/B _12633_/B _12606_/C VGND VGND VPWR VPWR _12607_/A sky130_fd_sc_hd__and3b_1
XFILLER_9_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13586_ _14108_/CLK hold249/X VGND VGND VPWR VPWR _13586_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10798_ _10798_/A VGND VGND VPWR VPWR _13061_/D sky130_fd_sc_hd__clkbuf_1
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12537_ _11317_/X _14714_/Q _12543_/S VGND VGND VPWR VPWR _12538_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12468_ _14665_/Q _12007_/A _12472_/S VGND VGND VPWR VPWR _12469_/A sky130_fd_sc_hd__mux2_1
X_14207_ _14209_/CLK _14207_/D VGND VGND VPWR VPWR _14207_/Q sky130_fd_sc_hd__dfxtp_1
X_11419_ _13732_/Q _11427_/B VGND VGND VPWR VPWR _11420_/A sky130_fd_sc_hd__and2_1
X_12399_ _12399_/A VGND VGND VPWR VPWR _14626_/D sky130_fd_sc_hd__clkbuf_1
X_14138_ _14716_/CLK _14138_/D VGND VGND VPWR VPWR hold412/A sky130_fd_sc_hd__dfxtp_1
XFILLER_113_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14069_ _14510_/CLK _14069_/D VGND VGND VPWR VPWR _14069_/Q sky130_fd_sc_hd__dfxtp_1
X_06960_ _07988_/B VGND VGND VPWR VPWR _08002_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_140_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _14667_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05911_ _05911_/A _05911_/B VGND VGND VPWR VPWR _06091_/A sky130_fd_sc_hd__nor2_1
XFILLER_95_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06891_ _06954_/A VGND VGND VPWR VPWR _07989_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_66_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08630_ _08630_/A _08630_/B _08630_/C _08630_/D VGND VGND VPWR VPWR _08630_/Y sky130_fd_sc_hd__nand4_1
XFILLER_54_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08561_ _08561_/A _08561_/B VGND VGND VPWR VPWR _08561_/Y sky130_fd_sc_hd__xnor2_1
X_07512_ _07532_/A _07510_/B _07503_/A VGND VGND VPWR VPWR _07519_/A sky130_fd_sc_hd__o21a_1
X_08492_ _09367_/B _08490_/B _08489_/X VGND VGND VPWR VPWR _08497_/B sky130_fd_sc_hd__o21bai_1
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07443_ _07443_/A _07443_/B VGND VGND VPWR VPWR _07454_/B sky130_fd_sc_hd__or2_1
XFILLER_11_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07374_ _07374_/A _07374_/B VGND VGND VPWR VPWR _07375_/C sky130_fd_sc_hd__and2_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09113_ _13527_/Q _09113_/B VGND VGND VPWR VPWR _09114_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06325_ _14404_/Q _14396_/Q _10197_/A VGND VGND VPWR VPWR _06325_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09044_ _09044_/A VGND VGND VPWR VPWR _12757_/D sky130_fd_sc_hd__clkbuf_1
X_06256_ _13954_/Q _13946_/Q _06256_/S VGND VGND VPWR VPWR _06256_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold420 hold420/A VGND VGND VPWR VPWR hold420/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06187_ _14417_/Q _14415_/Q _14426_/Q VGND VGND VPWR VPWR _06187_/X sky130_fd_sc_hd__mux2_1
Xhold431 hold431/A VGND VGND VPWR VPWR hold431/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_150_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold442 hold442/A VGND VGND VPWR VPWR hold442/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_145_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold453 hold453/A VGND VGND VPWR VPWR hold453/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold464 input18/X VGND VGND VPWR VPWR hold464/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold475 hold475/A VGND VGND VPWR VPWR hold475/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold486 hold486/A VGND VGND VPWR VPWR hold486/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_143_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold497 hold497/A VGND VGND VPWR VPWR hold497/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_09946_ _13497_/Q _13686_/Q _09946_/S VGND VGND VPWR VPWR _09947_/A sky130_fd_sc_hd__mux2_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _13691_/Q _09881_/D _09855_/X VGND VGND VPWR VPWR _09878_/B sky130_fd_sc_hd__o21ai_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08828_ _08828_/A _08953_/A VGND VGND VPWR VPWR _08847_/A sky130_fd_sc_hd__nand2_1
XFILLER_161_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08759_ _13461_/Q _09555_/B VGND VGND VPWR VPWR _08767_/A sky130_fd_sc_hd__nand2_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _13558_/Q _11772_/B VGND VGND VPWR VPWR _11771_/A sky130_fd_sc_hd__and2_1
XFILLER_72_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _10721_/A VGND VGND VPWR VPWR _12938_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _13702_/CLK _13440_/D repeater56/X VGND VGND VPWR VPWR _13440_/Q sky130_fd_sc_hd__dfrtp_1
X_10652_ _10652_/A VGND VGND VPWR VPWR _12679_/D sky130_fd_sc_hd__clkbuf_1
X_13371_ _13372_/CLK _13371_/D repeater57/X VGND VGND VPWR VPWR _13371_/Q sky130_fd_sc_hd__dfrtp_1
X_10583_ _10583_/A VGND VGND VPWR VPWR _13168_/D sky130_fd_sc_hd__clkbuf_1
X_12322_ _14576_/Q _12010_/X _12324_/S VGND VGND VPWR VPWR _12323_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12253_ _11317_/X _14542_/Q _12259_/S VGND VGND VPWR VPWR _12254_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11204_ _11159_/X _11201_/Y _11203_/Y _11166_/X VGND VGND VPWR VPWR _11205_/B sky130_fd_sc_hd__a211o_1
X_12184_ _12184_/A VGND VGND VPWR VPWR _14503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11135_ _13331_/Q _11079_/X _11128_/X _11134_/Y VGND VGND VPWR VPWR _13331_/D sky130_fd_sc_hd__o22a_1
XFILLER_150_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11066_ _11208_/A VGND VGND VPWR VPWR _11066_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10017_ _10052_/A _13913_/Q VGND VGND VPWR VPWR _10056_/A sky130_fd_sc_hd__xnor2_2
XFILLER_91_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11968_ _14699_/Q VGND VGND VPWR VPWR _11968_/X sky130_fd_sc_hd__clkbuf_2
X_13707_ _14645_/CLK _13707_/D VGND VGND VPWR VPWR _13707_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10919_ _14295_/Q _14465_/Q _14221_/Q _14051_/Q _10914_/X _12643_/A VGND VGND VPWR
+ VPWR _10919_/X sky130_fd_sc_hd__mux4_1
X_14687_ _14687_/CLK hold90/X VGND VGND VPWR VPWR _14687_/Q sky130_fd_sc_hd__dfxtp_2
X_11899_ _14257_/Q _11446_/X _11907_/S VGND VGND VPWR VPWR _11900_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13638_ _13653_/CLK hold337/X VGND VGND VPWR VPWR _13638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13569_ _14098_/CLK hold165/X VGND VGND VPWR VPWR _13569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06110_ _13783_/Q _13784_/Q _13785_/Q _13786_/Q VGND VGND VPWR VPWR _06110_/X sky130_fd_sc_hd__or4_1
XFILLER_8_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07090_ hold425/A _13706_/Q _07141_/B hold154/A VGND VGND VPWR VPWR _07093_/B sky130_fd_sc_hd__and4_1
XFILLER_146_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06041_ _06041_/A _06041_/B VGND VGND VPWR VPWR _10601_/A sky130_fd_sc_hd__nor2_1
XFILLER_145_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09800_ _09787_/S _09700_/X _09701_/X _09836_/D VGND VGND VPWR VPWR _09802_/B sky130_fd_sc_hd__o211a_1
X_07992_ _07998_/A _07992_/B _07992_/C VGND VGND VPWR VPWR _07992_/Y sky130_fd_sc_hd__nand3_1
XFILLER_113_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06943_ _06936_/A _06934_/X _06950_/A _06935_/A VGND VGND VPWR VPWR _06943_/X sky130_fd_sc_hd__a211o_1
X_09731_ _09731_/A VGND VGND VPWR VPWR _09836_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09662_ _14220_/Q _14218_/Q _14216_/Q _14214_/Q _09688_/S _13710_/Q VGND VGND VPWR
+ VPWR _09768_/B sky130_fd_sc_hd__mux4_2
X_06874_ _06976_/A VGND VGND VPWR VPWR _06874_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_82_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08613_ _13445_/Q _09438_/B _08620_/A _08601_/B VGND VGND VPWR VPWR _08614_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09593_ _09593_/A VGND VGND VPWR VPWR _12811_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08544_ _08544_/A VGND VGND VPWR VPWR _08544_/X sky130_fd_sc_hd__buf_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08475_ _08434_/Y _08595_/B _08474_/X _08431_/X VGND VGND VPWR VPWR _08490_/B sky130_fd_sc_hd__a22oi_4
X_07426_ _07455_/A _09163_/B VGND VGND VPWR VPWR _07426_/X sky130_fd_sc_hd__and2_1
XFILLER_50_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07357_ _07367_/A _07338_/X VGND VGND VPWR VPWR _07358_/B sky130_fd_sc_hd__or2b_1
XFILLER_164_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06308_ _06308_/A VGND VGND VPWR VPWR _14188_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07288_ _07350_/A _09099_/B VGND VGND VPWR VPWR _09098_/B sky130_fd_sc_hd__nor2_1
XFILLER_40_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09027_ _13214_/Q _13443_/Q _09029_/S VGND VGND VPWR VPWR _09028_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06239_ _14090_/Q _12036_/B VGND VGND VPWR VPWR _06240_/A sky130_fd_sc_hd__and2_1
XFILLER_151_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold250 hold250/A VGND VGND VPWR VPWR hold250/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold261 hold261/A VGND VGND VPWR VPWR hold261/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold272 hold272/A VGND VGND VPWR VPWR hold272/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_160_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold283 hold283/A VGND VGND VPWR VPWR hold283/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold294 hold294/A VGND VGND VPWR VPWR hold294/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09929_ _13489_/Q _13678_/Q _09935_/S VGND VGND VPWR VPWR _09930_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12940_ _13274_/CLK _12940_/D VGND VGND VPWR VPWR hold170/A sky130_fd_sc_hd__dfxtp_1
XFILLER_105_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _13698_/CLK _12871_/D VGND VGND VPWR VPWR hold155/A sky130_fd_sc_hd__dfxtp_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _14610_/CLK _14610_/D VGND VGND VPWR VPWR _14610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _13581_/Q _11828_/B VGND VGND VPWR VPWR _11823_/A sky130_fd_sc_hd__and2_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _11753_/A VGND VGND VPWR VPWR _14067_/D sky130_fd_sc_hd__clkbuf_1
X_14541_ _14713_/CLK _14541_/D VGND VGND VPWR VPWR _14541_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _10704_/A VGND VGND VPWR VPWR _12930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14472_ _14495_/CLK _14472_/D VGND VGND VPWR VPWR _14472_/Q sky130_fd_sc_hd__dfxtp_1
X_11684_ _11684_/A VGND VGND VPWR VPWR _14024_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10635_ _13814_/Q _10635_/B VGND VGND VPWR VPWR _13779_/D sky130_fd_sc_hd__xor2_1
X_13423_ _13423_/CLK hold477/X VGND VGND VPWR VPWR _13423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13354_ _13657_/CLK _13354_/D hold1/X VGND VGND VPWR VPWR _13354_/Q sky130_fd_sc_hd__dfrtp_1
X_10566_ _10567_/A _10573_/C VGND VGND VPWR VPWR _10566_/X sky130_fd_sc_hd__or2_1
XFILLER_6_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12305_ _14568_/Q _11984_/X _12313_/S VGND VGND VPWR VPWR _12306_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13285_ _13525_/CLK hold257/X VGND VGND VPWR VPWR _13285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10497_ _10498_/A _10498_/B _10498_/C VGND VGND VPWR VPWR _10503_/B sky130_fd_sc_hd__a21o_1
XFILLER_108_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12236_ _12236_/A VGND VGND VPWR VPWR _14534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12167_ _12167_/A VGND VGND VPWR VPWR _14495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11118_ _11118_/A VGND VGND VPWR VPWR _11118_/Y sky130_fd_sc_hd__inv_2
X_12098_ _14465_/Q _11950_/X _12106_/S VGND VGND VPWR VPWR _12099_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11049_ _14264_/Q _14655_/Q _13762_/Q _14710_/Q _11020_/X _11021_/X VGND VGND VPWR
+ VPWR _11050_/B sky130_fd_sc_hd__mux4_1
XFILLER_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 data_i[15] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__buf_6
XFILLER_36_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06590_ _06590_/A _06590_/B VGND VGND VPWR VPWR _12896_/D sky130_fd_sc_hd__nor2_1
XFILLER_80_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14739_ _14746_/CLK _14739_/D VGND VGND VPWR VPWR _14739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08260_ _09116_/S VGND VGND VPWR VPWR _08338_/A sky130_fd_sc_hd__buf_2
XFILLER_60_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07211_ _07211_/A VGND VGND VPWR VPWR _13351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08191_ _13359_/Q _08180_/B _08190_/X VGND VGND VPWR VPWR _08191_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07142_ _07142_/A _07142_/B VGND VGND VPWR VPWR _07144_/A sky130_fd_sc_hd__nor2_1
X_07073_ _07073_/A _07073_/B VGND VGND VPWR VPWR _07075_/A sky130_fd_sc_hd__nor2_1
XFILLER_146_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06024_ _14687_/Q _14683_/Q _14684_/Q _14685_/Q VGND VGND VPWR VPWR _06025_/B sky130_fd_sc_hd__and4_1
XFILLER_105_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07975_ _07975_/A _07975_/B VGND VGND VPWR VPWR _07975_/Y sky130_fd_sc_hd__nor2_1
X_06926_ _13014_/Q _13015_/Q _13016_/Q _13017_/Q _07988_/B VGND VGND VPWR VPWR _06926_/X
+ sky130_fd_sc_hd__o41a_1
X_09714_ _09718_/A VGND VGND VPWR VPWR _09735_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09645_ _13418_/Q _13616_/Q _09653_/S VGND VGND VPWR VPWR _09646_/A sky130_fd_sc_hd__mux2_1
X_06857_ _06857_/A _06857_/B VGND VGND VPWR VPWR _06876_/A sky130_fd_sc_hd__or2_1
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ _13619_/Q _09576_/B VGND VGND VPWR VPWR _09577_/B sky130_fd_sc_hd__or2_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06788_ _06770_/A _06786_/B _06770_/C _06785_/B VGND VGND VPWR VPWR _07863_/C sky130_fd_sc_hd__a31o_2
XFILLER_35_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _08527_/A _08527_/B VGND VGND VPWR VPWR _08531_/A sky130_fd_sc_hd__or2_1
XFILLER_35_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08458_ _13435_/Q _09370_/B VGND VGND VPWR VPWR _08459_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07409_ _08157_/A _09153_/B _09153_/C VGND VGND VPWR VPWR _07409_/X sky130_fd_sc_hd__and3_1
X_08389_ _13091_/Q _13372_/Q _08395_/S VGND VGND VPWR VPWR _08390_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10420_ _10421_/A _10421_/B _10421_/C VGND VGND VPWR VPWR _10426_/B sky130_fd_sc_hd__o21a_1
X_10351_ _06502_/A _13120_/D _10350_/X VGND VGND VPWR VPWR _10352_/B sky130_fd_sc_hd__o21ai_1
XFILLER_152_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13070_ _14082_/CLK _13070_/D VGND VGND VPWR VPWR hold239/A sky130_fd_sc_hd__dfxtp_1
X_10282_ _14326_/Q _14324_/Q _14595_/Q VGND VGND VPWR VPWR _10282_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12021_ _12021_/A VGND VGND VPWR VPWR _14316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13972_ _13972_/CLK _13972_/D VGND VGND VPWR VPWR _13972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12923_ _13039_/CLK _12923_/D VGND VGND VPWR VPWR hold423/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12854_ _13727_/CLK _12854_/D VGND VGND VPWR VPWR hold314/A sky130_fd_sc_hd__dfxtp_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _11805_/A VGND VGND VPWR VPWR _14095_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _13303_/CLK _12785_/D VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__dfxtp_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14524_ _14557_/CLK _14524_/D VGND VGND VPWR VPWR _14524_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ _11310_/X _14060_/Q _11736_/S VGND VGND VPWR VPWR _11737_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14455_ _14717_/CLK _14455_/D VGND VGND VPWR VPWR _14455_/Q sky130_fd_sc_hd__dfxtp_1
X_11667_ _14017_/Q _11462_/X _11667_/S VGND VGND VPWR VPWR _11668_/A sky130_fd_sc_hd__mux2_1
X_13406_ _13604_/CLK hold485/X VGND VGND VPWR VPWR _13406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10618_ _14196_/Q _14169_/Q _10617_/A VGND VGND VPWR VPWR _10618_/X sky130_fd_sc_hd__or3b_1
X_11598_ _14736_/Q VGND VGND VPWR VPWR _11655_/A sky130_fd_sc_hd__clkbuf_2
X_14386_ _14413_/CLK _14386_/D VGND VGND VPWR VPWR _14386_/Q sky130_fd_sc_hd__dfxtp_1
X_10549_ _10549_/A _10549_/B _10549_/C VGND VGND VPWR VPWR _10550_/B sky130_fd_sc_hd__and3_1
X_13337_ _14722_/CLK _13337_/D VGND VGND VPWR VPWR _13337_/Q sky130_fd_sc_hd__dfxtp_4
X_14763__74 VGND VGND VPWR VPWR _14763__74/HI _12911_/D sky130_fd_sc_hd__conb_1
XFILLER_6_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13268_ _13273_/CLK _13268_/D repeater59/X VGND VGND VPWR VPWR _13268_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12219_ _14124_/Q _12220_/C _12218_/Y VGND VGND VPWR VPWR _14517_/D sky130_fd_sc_hd__a21oi_1
X_13199_ _14333_/CLK _13199_/D VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07760_ _07760_/A _07760_/B VGND VGND VPWR VPWR _07761_/A sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_2_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06711_ _06681_/A _06681_/B _06698_/Y _06696_/Y VGND VGND VPWR VPWR _06712_/C sky130_fd_sc_hd__o211a_1
XFILLER_65_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07691_ _13112_/Q _07723_/C _07745_/B _13111_/Q VGND VGND VPWR VPWR _07693_/A sky130_fd_sc_hd__a22oi_1
XFILLER_37_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09430_ _08517_/X _08592_/X _09428_/Y _09429_/X VGND VGND VPWR VPWR _13598_/D sky130_fd_sc_hd__a22o_1
X_06642_ _13034_/Q VGND VGND VPWR VPWR _06643_/A sky130_fd_sc_hd__inv_2
XFILLER_53_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09361_ _13316_/Q _13554_/Q _10822_/A VGND VGND VPWR VPWR _09362_/A sky130_fd_sc_hd__mux2_1
X_06573_ _06567_/Y _06560_/B _06569_/A _06572_/X VGND VGND VPWR VPWR _06584_/C sky130_fd_sc_hd__a31o_1
XFILLER_33_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08312_ _08312_/A VGND VGND VPWR VPWR _08312_/Y sky130_fd_sc_hd__inv_2
X_09292_ _09290_/Y _09291_/X _07499_/A VGND VGND VPWR VPWR _13554_/D sky130_fd_sc_hd__o21bai_1
XFILLER_21_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_12 hold42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 input28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08243_ _13365_/Q _08243_/B VGND VGND VPWR VPWR _08256_/A sky130_fd_sc_hd__or2_1
XANTENNA_34 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_45 _13322_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 input8/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 _13548_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 _12004_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08174_ _13477_/Q _14011_/Q _08197_/A VGND VGND VPWR VPWR _08262_/B sky130_fd_sc_hd__mux2_1
XANTENNA_89 _13085_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07125_ _07151_/A _07123_/Y _07093_/B _07107_/C VGND VGND VPWR VPWR _07128_/B sky130_fd_sc_hd__a211o_1
XFILLER_161_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07056_ _07034_/Y _07055_/Y _10647_/A VGND VGND VPWR VPWR _07057_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06007_ _13559_/Q _13560_/Q _13561_/Q _13562_/Q VGND VGND VPWR VPWR _06007_/X sky130_fd_sc_hd__and4_1
XFILLER_133_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07958_ _07948_/A _07952_/X _07972_/B VGND VGND VPWR VPWR _07958_/X sky130_fd_sc_hd__a21o_1
XFILLER_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06909_ _06909_/A _06904_/B VGND VGND VPWR VPWR _06914_/B sky130_fd_sc_hd__or2b_1
X_07889_ _13264_/Q _07889_/B VGND VGND VPWR VPWR _07890_/B sky130_fd_sc_hd__or2_1
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09628_ _09628_/A VGND VGND VPWR VPWR _12827_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09559_ _09559_/A _09559_/B VGND VGND VPWR VPWR _09559_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12570_ _14742_/Q VGND VGND VPWR VPWR _12570_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11521_ _11521_/A VGND VGND VPWR VPWR _13841_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14240_ _14510_/CLK _14240_/D VGND VGND VPWR VPWR _14240_/Q sky130_fd_sc_hd__dfxtp_1
X_11452_ _11452_/A VGND VGND VPWR VPWR _13819_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10403_ _10386_/A _13519_/Q _13520_/Q _13516_/Q VGND VGND VPWR VPWR _10403_/X sky130_fd_sc_hd__a22o_1
X_14171_ _14196_/CLK _14171_/D VGND VGND VPWR VPWR _14171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11383_ _11383_/A VGND VGND VPWR VPWR _13785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13122_ _13666_/CLK _14634_/Q VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__dfxtp_1
XFILLER_3_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10334_ _10334_/A _10334_/B VGND VGND VPWR VPWR _13172_/D sky130_fd_sc_hd__xnor2_1
XFILLER_152_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ _13565_/CLK _13053_/D VGND VGND VPWR VPWR hold417/A sky130_fd_sc_hd__dfxtp_1
X_10265_ _10265_/A VGND VGND VPWR VPWR _14354_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12004_ _12004_/A VGND VGND VPWR VPWR _12004_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10196_ _14397_/Q _14389_/Q _10197_/A VGND VGND VPWR VPWR _10626_/C sky130_fd_sc_hd__mux2_1
XFILLER_66_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13955_ _13972_/CLK _13955_/D VGND VGND VPWR VPWR _13955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12906_ _13280_/CLK _12906_/D repeater59/X VGND VGND VPWR VPWR _12906_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13886_ _14210_/CLK hold316/X VGND VGND VPWR VPWR _13886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _14656_/CLK _12837_/D VGND VGND VPWR VPWR hold328/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _13855_/CLK _12768_/D VGND VGND VPWR VPWR hold435/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _14579_/CLK _14507_/D VGND VGND VPWR VPWR _14507_/Q sky130_fd_sc_hd__dfxtp_1
X_11719_ _11285_/X _14052_/Q _11725_/S VGND VGND VPWR VPWR _11720_/A sky130_fd_sc_hd__mux2_1
X_12699_ _13027_/CLK _12699_/D VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__dfxtp_1
X_14438_ _14439_/CLK _14438_/D VGND VGND VPWR VPWR _14438_/Q sky130_fd_sc_hd__dfxtp_1
Xinput10 data_i[18] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__buf_2
XFILLER_163_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput21 data_i[4] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__buf_2
X_14369_ _14425_/CLK _14369_/D VGND VGND VPWR VPWR _14369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08930_ _08930_/A _08930_/B VGND VGND VPWR VPWR _08932_/A sky130_fd_sc_hd__nor2_1
XFILLER_112_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08861_ _08861_/A _08861_/B VGND VGND VPWR VPWR _08863_/A sky130_fd_sc_hd__nor2_1
XFILLER_97_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07812_ _13252_/Q _07807_/B _07805_/X _07806_/A VGND VGND VPWR VPWR _07815_/A sky130_fd_sc_hd__a31o_1
XFILLER_69_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08792_ _08784_/X _08790_/X _08791_/Y _08764_/X VGND VGND VPWR VPWR _13465_/D sky130_fd_sc_hd__a31o_1
X_07743_ _07772_/A _07772_/B VGND VGND VPWR VPWR _07745_/C sky130_fd_sc_hd__and2_1
XFILLER_84_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07674_ _07675_/A _07675_/B _07675_/C VGND VGND VPWR VPWR _07689_/B sky130_fd_sc_hd__o21a_1
XFILLER_37_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06625_ _12907_/Q _06620_/X _06624_/Y VGND VGND VPWR VPWR _12907_/D sky130_fd_sc_hd__a21oi_1
X_09413_ _09413_/A VGND VGND VPWR VPWR _13596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09344_ _09344_/A VGND VGND VPWR VPWR _12798_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06556_ _12890_/Q _06556_/B VGND VGND VPWR VPWR _06557_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09275_ _09273_/Y _09274_/X _07499_/A VGND VGND VPWR VPWR _13551_/D sky130_fd_sc_hd__o21bai_1
X_06487_ _06493_/B _06499_/A VGND VGND VPWR VPWR _06490_/A sky130_fd_sc_hd__nor2_1
XFILLER_138_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08226_ _09125_/A _08226_/B VGND VGND VPWR VPWR _08226_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08157_ _08157_/A VGND VGND VPWR VPWR _08157_/X sky130_fd_sc_hd__buf_4
XFILLER_146_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07108_ _14630_/Q VGND VGND VPWR VPWR _07163_/B sky130_fd_sc_hd__clkbuf_2
X_08088_ _08088_/A VGND VGND VPWR VPWR _12703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07039_ _13707_/Q VGND VGND VPWR VPWR _07165_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_164_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10050_ _13805_/Q _13789_/Q _10050_/S VGND VGND VPWR VPWR _10051_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13740_ _13811_/CLK hold388/X VGND VGND VPWR VPWR _13740_/Q sky130_fd_sc_hd__dfxtp_1
X_10952_ _10952_/A _10925_/X VGND VGND VPWR VPWR _10952_/X sky130_fd_sc_hd__or2b_1
XFILLER_73_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13671_ _13673_/CLK _13671_/D repeater56/X VGND VGND VPWR VPWR _13671_/Q sky130_fd_sc_hd__dfrtp_1
X_10883_ _13158_/Q _10885_/B VGND VGND VPWR VPWR _10884_/A sky130_fd_sc_hd__and2_1
X_12622_ _14733_/Q _12616_/B _12621_/X _12617_/X VGND VGND VPWR VPWR _14738_/D sky130_fd_sc_hd__o211a_1
X_12553_ _12553_/A VGND VGND VPWR VPWR _14721_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11504_ _12007_/A VGND VGND VPWR VPWR _11504_/X sky130_fd_sc_hd__clkbuf_2
X_12484_ _12484_/A _12484_/B input9/X VGND VGND VPWR VPWR _12485_/A sky130_fd_sc_hd__and3_1
XFILLER_156_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14223_ _14535_/CLK _14223_/D VGND VGND VPWR VPWR _14223_/Q sky130_fd_sc_hd__dfxtp_1
X_11435_ _11435_/A VGND VGND VPWR VPWR _13808_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14154_ _14294_/CLK hold383/X VGND VGND VPWR VPWR _14154_/Q sky130_fd_sc_hd__dfxtp_1
X_11366_ _13776_/Q _11365_/X _11376_/S VGND VGND VPWR VPWR _11367_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13105_ _13294_/CLK hold245/X VGND VGND VPWR VPWR _13105_/Q sky130_fd_sc_hd__dfxtp_1
X_10317_ _10317_/A _10317_/B VGND VGND VPWR VPWR _13476_/D sky130_fd_sc_hd__xnor2_1
XFILLER_140_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11297_ _14699_/Q VGND VGND VPWR VPWR _11297_/X sky130_fd_sc_hd__buf_2
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14085_ _14397_/CLK _14085_/D VGND VGND VPWR VPWR _14085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ _14527_/D _10247_/X _14556_/D VGND VGND VPWR VPWR _10248_/X sky130_fd_sc_hd__mux2_1
X_13036_ _13353_/CLK _13036_/D VGND VGND VPWR VPWR _13036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10179_ _10172_/X _14140_/D _10179_/S VGND VGND VPWR VPWR _10179_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13938_ _13972_/CLK _13938_/D VGND VGND VPWR VPWR _13938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13869_ _14075_/CLK _13869_/D VGND VGND VPWR VPWR _13869_/Q sky130_fd_sc_hd__dfxtp_1
X_06410_ _14437_/Q _14435_/Q _06425_/S VGND VGND VPWR VPWR _06410_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07390_ _07401_/A _07401_/B VGND VGND VPWR VPWR _07395_/A sky130_fd_sc_hd__xor2_2
XFILLER_148_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06341_ _14107_/Q _14091_/Q _06341_/S VGND VGND VPWR VPWR _06342_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09060_ _13228_/Q _13457_/Q _09064_/S VGND VGND VPWR VPWR _09061_/A sky130_fd_sc_hd__mux2_1
X_06272_ _06272_/A VGND VGND VPWR VPWR _13954_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08011_ _06793_/A _08009_/Y _08010_/X _06930_/X VGND VGND VPWR VPWR _13281_/D sky130_fd_sc_hd__a31o_1
XFILLER_163_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09962_ _13504_/Q _13693_/Q _09968_/S VGND VGND VPWR VPWR _09963_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08913_ _08939_/A _08911_/Y _08881_/B _08895_/C VGND VGND VPWR VPWR _08916_/B sky130_fd_sc_hd__a211o_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _09893_/A _09893_/B VGND VGND VPWR VPWR _09894_/C sky130_fd_sc_hd__nand2_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08844_ _08822_/Y _08843_/Y _11268_/A VGND VGND VPWR VPWR _08845_/A sky130_fd_sc_hd__mux2_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05987_ _05987_/A _05987_/B _05987_/C VGND VGND VPWR VPWR _05994_/A sky130_fd_sc_hd__nor3_1
X_08775_ _08775_/A _08775_/B VGND VGND VPWR VPWR _08786_/B sky130_fd_sc_hd__or2_1
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07726_ _07726_/A _07726_/B VGND VGND VPWR VPWR _07753_/B sky130_fd_sc_hd__xnor2_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07657_ _07657_/A _07657_/B VGND VGND VPWR VPWR _07659_/C sky130_fd_sc_hd__xor2_1
XFILLER_41_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06608_ _12900_/Q _12901_/Q _06607_/D _12902_/Q VGND VGND VPWR VPWR _06609_/C sky130_fd_sc_hd__a31o_1
X_07588_ _07585_/Y _07586_/X _07581_/A _07587_/Y VGND VGND VPWR VPWR _07588_/X sky130_fd_sc_hd__a211o_1
X_09327_ _09327_/A VGND VGND VPWR VPWR _12790_/D sky130_fd_sc_hd__clkbuf_1
X_06539_ _12910_/Q VGND VGND VPWR VPWR _06599_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09258_ _13549_/Q _09258_/B VGND VGND VPWR VPWR _09259_/B sky130_fd_sc_hd__or2_1
XFILLER_138_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08209_ _13362_/Q _08209_/B _08250_/C VGND VGND VPWR VPWR _08211_/A sky130_fd_sc_hd__and3_1
X_09189_ _09189_/A _09189_/B VGND VGND VPWR VPWR _09190_/B sky130_fd_sc_hd__nor2_1
XFILLER_107_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11220_ _13337_/Q _11150_/X _11213_/X _11219_/Y VGND VGND VPWR VPWR _13337_/D sky130_fd_sc_hd__o22a_1
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11151_ _14310_/Q _14480_/Q _14236_/Q _14066_/Q _11137_/X _11138_/X VGND VGND VPWR
+ VPWR _11151_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10102_ _10139_/A _14144_/Q VGND VGND VPWR VPWR _10103_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11082_ _11153_/A VGND VGND VPWR VPWR _11082_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10033_ _10033_/A VGND VGND VPWR VPWR _13970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11984_ _14515_/Q VGND VGND VPWR VPWR _11984_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13723_ _13727_/CLK hold83/X VGND VGND VPWR VPWR _13723_/Q sky130_fd_sc_hd__dfxtp_1
X_10935_ _14746_/Q VGND VGND VPWR VPWR _11153_/A sky130_fd_sc_hd__buf_4
XFILLER_16_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13654_ _14693_/CLK hold48/X VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10866_ _13150_/Q _10874_/B VGND VGND VPWR VPWR _10867_/A sky130_fd_sc_hd__and2_1
XFILLER_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12605_ _12616_/A _14730_/Q _12623_/B _14732_/Q VGND VGND VPWR VPWR _12606_/C sky130_fd_sc_hd__a31o_1
XFILLER_31_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13585_ _14108_/CLK hold347/X VGND VGND VPWR VPWR _13585_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10797_ _13019_/Q _10801_/B VGND VGND VPWR VPWR _10798_/A sky130_fd_sc_hd__and2_1
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12536_ _12536_/A VGND VGND VPWR VPWR _14713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12467_ _12467_/A VGND VGND VPWR VPWR _14664_/D sky130_fd_sc_hd__clkbuf_1
X_14206_ _14208_/CLK _14206_/D VGND VGND VPWR VPWR _14206_/Q sky130_fd_sc_hd__dfxtp_1
X_11418_ _11429_/A VGND VGND VPWR VPWR _11427_/B sky130_fd_sc_hd__clkbuf_1
X_12398_ input12/X _12402_/B _12400_/C VGND VGND VPWR VPWR _12399_/A sky130_fd_sc_hd__and3_1
XFILLER_153_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14137_ _14159_/CLK _14137_/D VGND VGND VPWR VPWR hold292/A sky130_fd_sc_hd__dfxtp_1
X_11349_ _13773_/Q _11348_/X _11355_/S VGND VGND VPWR VPWR _11350_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14068_ _14510_/CLK _14068_/D VGND VGND VPWR VPWR _14068_/Q sky130_fd_sc_hd__dfxtp_1
X_13019_ _13570_/CLK _13019_/D repeater59/X VGND VGND VPWR VPWR _13019_/Q sky130_fd_sc_hd__dfrtp_1
X_05910_ _13800_/Q _13801_/Q _05910_/C _05910_/D VGND VGND VPWR VPWR _05911_/B sky130_fd_sc_hd__and4_1
X_06890_ _07968_/B VGND VGND VPWR VPWR _06954_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08560_ _08572_/A _08539_/X VGND VGND VPWR VPWR _08561_/B sky130_fd_sc_hd__or2b_1
XFILLER_35_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07511_ _07495_/X _07509_/X _07510_/Y _07499_/X VGND VGND VPWR VPWR _13151_/D sky130_fd_sc_hd__a31o_1
X_08491_ _08582_/A VGND VGND VPWR VPWR _08567_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_07442_ _07442_/A _07442_/B VGND VGND VPWR VPWR _07443_/B sky130_fd_sc_hd__or2_1
X_07373_ _07387_/A _07372_/X _07363_/B VGND VGND VPWR VPWR _07374_/B sky130_fd_sc_hd__o21a_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06324_ _06324_/A _06324_/B VGND VGND VPWR VPWR _06324_/Y sky130_fd_sc_hd__nand2_1
X_09112_ _13528_/Q _09112_/B VGND VGND VPWR VPWR _09134_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09043_ _13221_/Q _13450_/Q _09051_/S VGND VGND VPWR VPWR _09044_/A sky130_fd_sc_hd__mux2_1
X_06255_ _06255_/A VGND VGND VPWR VPWR _14412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold410 hold410/A VGND VGND VPWR VPWR hold410/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06186_ _14418_/Q _14416_/Q _14426_/Q VGND VGND VPWR VPWR _06186_/X sky130_fd_sc_hd__mux2_1
Xhold421 hold421/A VGND VGND VPWR VPWR hold421/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold432 hold432/A VGND VGND VPWR VPWR hold432/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold443 hold443/A VGND VGND VPWR VPWR hold443/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_145_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold454 hold454/A VGND VGND VPWR VPWR hold454/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold465 hold465/A VGND VGND VPWR VPWR hold465/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold476 hold476/A VGND VGND VPWR VPWR hold476/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold487 hold487/A VGND VGND VPWR VPWR hold487/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold498 hold498/A VGND VGND VPWR VPWR hold498/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09945_ _09945_/A VGND VGND VPWR VPWR _12859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09876_ _13691_/Q _09881_/D VGND VGND VPWR VPWR _09878_/A sky130_fd_sc_hd__and2_1
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _13518_/D VGND VGND VPWR VPWR _08953_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _08758_/A _08758_/B VGND VGND VPWR VPWR _08763_/C sky130_fd_sc_hd__nand2_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _07680_/A _07680_/B _07708_/Y VGND VGND VPWR VPWR _07710_/C sky130_fd_sc_hd__o21ai_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _08714_/A _08689_/B VGND VGND VPWR VPWR _08689_/X sky130_fd_sc_hd__and2b_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10720_ _12895_/Q _10720_/B VGND VGND VPWR VPWR _10721_/A sky130_fd_sc_hd__and2_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10651_ _13622_/Q _11529_/B VGND VGND VPWR VPWR _10652_/A sky130_fd_sc_hd__and2_1
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13370_ _13555_/CLK _13370_/D repeater57/X VGND VGND VPWR VPWR _13370_/Q sky130_fd_sc_hd__dfrtp_1
X_10582_ hold519/A hold507/X VGND VGND VPWR VPWR _10583_/A sky130_fd_sc_hd__or2_1
X_12321_ _12321_/A VGND VGND VPWR VPWR _14575_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12252_ _12252_/A VGND VGND VPWR VPWR _14541_/D sky130_fd_sc_hd__clkbuf_1
X_11203_ _11240_/A _11203_/B VGND VGND VPWR VPWR _11203_/Y sky130_fd_sc_hd__nor2_1
X_12183_ _14503_/Q _11997_/X _12183_/S VGND VGND VPWR VPWR _12184_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11134_ _11179_/A _11134_/B VGND VGND VPWR VPWR _11134_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11065_ _11262_/A VGND VGND VPWR VPWR _11065_/X sky130_fd_sc_hd__buf_2
XFILLER_1_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10016_ _10016_/A VGND VGND VPWR VPWR _14050_/D sky130_fd_sc_hd__inv_2
XFILLER_37_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11967_ _11967_/A VGND VGND VPWR VPWR _14299_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13706_ _14645_/CLK _13706_/D VGND VGND VPWR VPWR _13706_/Q sky130_fd_sc_hd__dfxtp_1
X_10918_ _10918_/A VGND VGND VPWR VPWR _12643_/A sky130_fd_sc_hd__buf_2
X_14686_ _14688_/CLK hold336/X VGND VGND VPWR VPWR _14686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11898_ _11948_/S VGND VGND VPWR VPWR _11907_/S sky130_fd_sc_hd__buf_2
XFILLER_20_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13637_ _13653_/CLK hold489/X VGND VGND VPWR VPWR _13637_/Q sky130_fd_sc_hd__dfxtp_1
X_10849_ _10849_/A VGND VGND VPWR VPWR _13184_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13568_ _13574_/CLK hold21/X VGND VGND VPWR VPWR _13568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12519_ _11291_/X _14706_/Q _12521_/S VGND VGND VPWR VPWR _12520_/A sky130_fd_sc_hd__mux2_1
X_13499_ _13700_/CLK hold202/X VGND VGND VPWR VPWR _13499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06040_ input20/X input21/X input22/X _06371_/B VGND VGND VPWR VPWR _06041_/B sky130_fd_sc_hd__o31a_1
XFILLER_114_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07991_ _07992_/B _07992_/C _07998_/A VGND VGND VPWR VPWR _07995_/B sky130_fd_sc_hd__a21o_1
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_7_0_clk clkbuf_4_7_0_clk/A VGND VGND VPWR VPWR clkbuf_4_7_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09730_ _09730_/A VGND VGND VPWR VPWR _13671_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06942_ _06948_/B VGND VGND VPWR VPWR _06942_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09661_ _13709_/Q VGND VGND VPWR VPWR _09688_/S sky130_fd_sc_hd__clkbuf_2
X_06873_ _07861_/S VGND VGND VPWR VPWR _06976_/A sky130_fd_sc_hd__buf_2
XFILLER_55_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08612_ _08620_/B _08620_/C VGND VGND VPWR VPWR _08614_/A sky130_fd_sc_hd__or2_1
XFILLER_54_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09592_ _13394_/Q _13592_/Q _09598_/S VGND VGND VPWR VPWR _09593_/A sky130_fd_sc_hd__mux2_2
XFILLER_36_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08543_ _08517_/X _09417_/B _08539_/X _08542_/Y VGND VGND VPWR VPWR _13441_/D sky130_fd_sc_hd__a22o_1
XFILLER_70_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08474_ _08645_/A _08471_/X _08473_/X VGND VGND VPWR VPWR _08474_/X sky130_fd_sc_hd__a21o_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07425_ _07425_/A _07425_/B _07425_/C _07425_/D VGND VGND VPWR VPWR _07425_/Y sky130_fd_sc_hd__nand4_1
XFILLER_11_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07356_ _13137_/Q _07356_/B VGND VGND VPWR VPWR _07367_/A sky130_fd_sc_hd__and2_1
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06307_ _13874_/Q _13858_/Q _06309_/S VGND VGND VPWR VPWR _06308_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07287_ _07261_/B _07284_/B _07283_/X VGND VGND VPWR VPWR _09099_/B sky130_fd_sc_hd__o21ba_1
XFILLER_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06238_ _06238_/A VGND VGND VPWR VPWR _14388_/D sky130_fd_sc_hd__clkbuf_1
X_09026_ _09026_/A VGND VGND VPWR VPWR _12749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06169_ _13858_/Q _11836_/B VGND VGND VPWR VPWR _06170_/A sky130_fd_sc_hd__and2_1
Xhold240 hold240/A VGND VGND VPWR VPWR hold240/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold251 hold251/A VGND VGND VPWR VPWR hold251/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold262 hold262/A VGND VGND VPWR VPWR hold262/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold273 hold273/A VGND VGND VPWR VPWR hold273/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold284 hold284/A VGND VGND VPWR VPWR hold284/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold295 hold295/A VGND VGND VPWR VPWR hold295/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09928_ _09928_/A VGND VGND VPWR VPWR _12851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09859_ _09873_/C VGND VGND VPWR VPWR _09870_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _13811_/CLK _12870_/D VGND VGND VPWR VPWR hold434/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _11821_/A VGND VGND VPWR VPWR _14102_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _14709_/CLK _14540_/D VGND VGND VPWR VPWR _14540_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _11337_/X _14067_/Q _11758_/S VGND VGND VPWR VPWR _11753_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _12887_/Q _10709_/B VGND VGND VPWR VPWR _10704_/A sky130_fd_sc_hd__and2_1
X_14471_ _14600_/CLK _14471_/D VGND VGND VPWR VPWR _14471_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _14024_/Q _11485_/X _11689_/S VGND VGND VPWR VPWR _11684_/A sky130_fd_sc_hd__mux2_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ _13617_/CLK hold109/X VGND VGND VPWR VPWR _13422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10634_ _10634_/A VGND VGND VPWR VPWR _14587_/D sky130_fd_sc_hd__clkinv_2
XFILLER_139_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13353_ _13353_/CLK _13353_/D VGND VGND VPWR VPWR _13353_/Q sky130_fd_sc_hd__dfxtp_1
X_10565_ _10565_/A _10560_/B VGND VGND VPWR VPWR _10570_/A sky130_fd_sc_hd__or2b_1
X_12304_ _12315_/A VGND VGND VPWR VPWR _12313_/S sky130_fd_sc_hd__buf_2
XFILLER_143_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13284_ _13294_/CLK _13284_/D hold1/X VGND VGND VPWR VPWR _13284_/Q sky130_fd_sc_hd__dfrtp_1
X_10496_ _10460_/A _10494_/X _10503_/A _10486_/B VGND VGND VPWR VPWR _10498_/C sky130_fd_sc_hd__a31oi_1
XFILLER_6_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12235_ _11291_/X _14534_/Q _12237_/S VGND VGND VPWR VPWR _12236_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12166_ _14495_/Q _11972_/X _12172_/S VGND VGND VPWR VPWR _12167_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11117_ _14608_/Q _14570_/Q _14501_/Q _14453_/Q _11115_/X _11116_/X VGND VGND VPWR
+ VPWR _11118_/A sky130_fd_sc_hd__mux4_1
X_12097_ _12147_/S VGND VGND VPWR VPWR _12106_/S sky130_fd_sc_hd__buf_2
XFILLER_1_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11048_ _11190_/A VGND VGND VPWR VPWR _11106_/A sky130_fd_sc_hd__clkbuf_2
Xinput8 data_i[16] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__buf_6
XFILLER_64_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12999_ _14647_/CLK _12999_/D hold1/X VGND VGND VPWR VPWR _12999_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_91_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14738_ _14746_/CLK _14738_/D VGND VGND VPWR VPWR _14738_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14669_ _14724_/CLK _14669_/D VGND VGND VPWR VPWR _14669_/Q sky130_fd_sc_hd__dfxtp_1
X_07210_ _07198_/Y _07209_/Y _07218_/S VGND VGND VPWR VPWR _07211_/A sky130_fd_sc_hd__mux2_1
X_08190_ _13358_/Q _08166_/B _08180_/B _13359_/Q VGND VGND VPWR VPWR _08190_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07141_ _07141_/A _07141_/B _07141_/C _07163_/B VGND VGND VPWR VPWR _07142_/B sky130_fd_sc_hd__and4_1
XFILLER_9_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07072_ _07072_/A _07072_/B VGND VGND VPWR VPWR _07073_/B sky130_fd_sc_hd__nor2_1
XFILLER_105_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06023_ _11772_/B VGND VGND VPWR VPWR _14380_/D sky130_fd_sc_hd__inv_2
XFILLER_114_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07974_ _13272_/Q _13273_/Q _13274_/Q _13275_/Q _07981_/B VGND VGND VPWR VPWR _07975_/B
+ sky130_fd_sc_hd__o41a_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09713_ _09713_/A VGND VGND VPWR VPWR _13670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06925_ _07989_/B VGND VGND VPWR VPWR _07988_/B sky130_fd_sc_hd__buf_2
XFILLER_95_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09644_ _09644_/A VGND VGND VPWR VPWR _09653_/S sky130_fd_sc_hd__clkbuf_2
X_06856_ _06857_/A _06858_/A _06857_/B VGND VGND VPWR VPWR _06856_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_27_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09575_ _13619_/Q _09576_/B VGND VGND VPWR VPWR _09577_/A sky130_fd_sc_hd__nand2_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06787_ _06813_/A VGND VGND VPWR VPWR _07863_/B sky130_fd_sc_hd__buf_2
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08526_ _13440_/Q _09401_/B VGND VGND VPWR VPWR _08527_/B sky130_fd_sc_hd__nor2_1
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08457_ _08457_/A _08457_/B VGND VGND VPWR VPWR _08459_/A sky130_fd_sc_hd__or2_1
XFILLER_51_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07408_ _07408_/A _07408_/B VGND VGND VPWR VPWR _07408_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_156_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08388_ _08388_/A VGND VGND VPWR VPWR _12726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07339_ _07473_/A VGND VGND VPWR VPWR _07341_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_137_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10350_ _06502_/A _13120_/D _10347_/A VGND VGND VPWR VPWR _10350_/X sky130_fd_sc_hd__a21bo_1
XFILLER_164_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09009_ _09655_/S VGND VGND VPWR VPWR _09018_/S sky130_fd_sc_hd__clkbuf_2
X_10281_ _10281_/A VGND VGND VPWR VPWR _12664_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12020_ _14316_/Q _12019_/X _12026_/S VGND VGND VPWR VPWR _12021_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13971_ _13978_/CLK _13971_/D VGND VGND VPWR VPWR _13971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12922_ _13039_/CLK _12922_/D VGND VGND VPWR VPWR hold252/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12853_ _13727_/CLK _12853_/D VGND VGND VPWR VPWR hold279/A sky130_fd_sc_hd__dfxtp_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _13573_/Q _11806_/B VGND VGND VPWR VPWR _11805_/A sky130_fd_sc_hd__and2_1
XFILLER_73_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _13294_/CLK _12784_/D VGND VGND VPWR VPWR hold103/A sky130_fd_sc_hd__dfxtp_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14523_ _14557_/CLK _14523_/D VGND VGND VPWR VPWR _14523_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _11735_/A VGND VGND VPWR VPWR _14059_/D sky130_fd_sc_hd__clkbuf_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14454_ _14610_/CLK _14454_/D VGND VGND VPWR VPWR _14454_/Q sky130_fd_sc_hd__dfxtp_1
X_11666_ _11666_/A VGND VGND VPWR VPWR _14016_/D sky130_fd_sc_hd__clkbuf_1
X_13405_ _13604_/CLK hold465/X VGND VGND VPWR VPWR _13405_/Q sky130_fd_sc_hd__dfxtp_1
X_10617_ _10617_/A _14177_/Q _14195_/Q VGND VGND VPWR VPWR _10617_/X sky130_fd_sc_hd__or3_1
X_14385_ _14413_/CLK hold125/X VGND VGND VPWR VPWR _14385_/Q sky130_fd_sc_hd__dfxtp_1
X_11597_ _11597_/A VGND VGND VPWR VPWR _13960_/D sky130_fd_sc_hd__inv_2
X_13336_ _14722_/CLK _13336_/D VGND VGND VPWR VPWR _13336_/Q sky130_fd_sc_hd__dfxtp_2
X_10548_ _10549_/A _10549_/B _10549_/C VGND VGND VPWR VPWR _10562_/A sky130_fd_sc_hd__a21oi_1
X_13267_ _13273_/CLK _13267_/D repeater59/X VGND VGND VPWR VPWR _13267_/Q sky130_fd_sc_hd__dfrtp_1
X_10479_ _10481_/A _10481_/B VGND VGND VPWR VPWR _14009_/D sky130_fd_sc_hd__xor2_1
X_12218_ _14124_/Q _12220_/C _12205_/X VGND VGND VPWR VPWR _12218_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_151_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13198_ _13617_/CLK _13198_/D VGND VGND VPWR VPWR hold447/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12149_ _12149_/A _11841_/A VGND VGND VPWR VPWR _12342_/B sky130_fd_sc_hd__or2b_2
XFILLER_111_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06710_ _13002_/Q _06710_/B VGND VGND VPWR VPWR _06712_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07690_ _14584_/Q VGND VGND VPWR VPWR _07745_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06641_ _07807_/B _06641_/B VGND VGND VPWR VPWR _12998_/D sky130_fd_sc_hd__xnor2_1
XFILLER_64_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09360_ _09360_/A VGND VGND VPWR VPWR _12805_/D sky130_fd_sc_hd__clkbuf_1
X_06572_ _06557_/A _06566_/A _06566_/B VGND VGND VPWR VPWR _06572_/X sky130_fd_sc_hd__o21ba_1
XFILLER_80_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08311_ _08314_/B _08317_/D VGND VGND VPWR VPWR _08312_/A sky130_fd_sc_hd__and2_1
XFILLER_61_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09291_ _09285_/A _09286_/X _09289_/Y _07396_/A VGND VGND VPWR VPWR _09291_/X sky130_fd_sc_hd__a31o_1
XFILLER_32_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_13 hold42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08242_ _13365_/Q _08243_/B VGND VGND VPWR VPWR _08244_/A sky130_fd_sc_hd__and2_1
XANTENNA_24 input29/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_35 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 _13326_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 input8/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 _13549_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08173_ _14009_/Q _14007_/Q _08197_/A VGND VGND VPWR VPWR _08173_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_79 _12016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07124_ _07093_/B _07107_/C _07151_/A _07123_/Y VGND VGND VPWR VPWR _07151_/B sky130_fd_sc_hd__o211ai_2
XFILLER_134_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07055_ _07156_/A _07055_/B VGND VGND VPWR VPWR _07055_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_118_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06006_ hold173/A _13564_/Q _06006_/C _06006_/D VGND VGND VPWR VPWR _06006_/X sky130_fd_sc_hd__and4_1
XFILLER_0_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07957_ _07957_/A _07957_/B VGND VGND VPWR VPWR _07972_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06908_ _06861_/X _06905_/X _06906_/Y _06907_/X VGND VGND VPWR VPWR _13015_/D sky130_fd_sc_hd__a31o_1
XFILLER_101_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07888_ _13264_/Q _07889_/B VGND VGND VPWR VPWR _07898_/A sky130_fd_sc_hd__nand2_1
XFILLER_44_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09627_ _13410_/Q _13608_/Q _09631_/S VGND VGND VPWR VPWR _09628_/A sky130_fd_sc_hd__mux2_1
X_06839_ _06846_/B _06837_/Y _06838_/X VGND VGND VPWR VPWR _13010_/D sky130_fd_sc_hd__a21o_1
XFILLER_55_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09558_ _08504_/X _09557_/Y _09493_/X VGND VGND VPWR VPWR _13616_/D sky130_fd_sc_hd__a21o_1
XFILLER_62_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08509_ _08521_/A _08509_/B VGND VGND VPWR VPWR _09394_/B sky130_fd_sc_hd__xor2_4
XFILLER_70_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09489_ _13606_/Q _09511_/B VGND VGND VPWR VPWR _09500_/A sky130_fd_sc_hd__nand2_1
X_11520_ _13841_/Q _11519_/X _11523_/S VGND VGND VPWR VPWR _11521_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11451_ _13819_/Q _11446_/X _11463_/S VGND VGND VPWR VPWR _11452_/A sky130_fd_sc_hd__mux2_1
X_10402_ _10423_/A _10429_/C VGND VGND VPWR VPWR _10431_/A sky130_fd_sc_hd__nand2_1
X_14170_ _14196_/CLK _14170_/D VGND VGND VPWR VPWR _14170_/Q sky130_fd_sc_hd__dfxtp_1
X_11382_ _13716_/Q _11382_/B VGND VGND VPWR VPWR _11383_/A sky130_fd_sc_hd__and2_1
XFILLER_152_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13121_ _13657_/CLK _13121_/D VGND VGND VPWR VPWR hold84/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10333_ _13108_/Q _13241_/D _10332_/X VGND VGND VPWR VPWR _10334_/B sky130_fd_sc_hd__o21ai_1
XFILLER_124_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13052_ _13565_/CLK _13052_/D VGND VGND VPWR VPWR hold365/A sky130_fd_sc_hd__dfxtp_1
X_10264_ _10260_/X _10263_/X _10269_/S VGND VGND VPWR VPWR _10265_/A sky130_fd_sc_hd__mux2_1
X_12003_ _12003_/A VGND VGND VPWR VPWR _14310_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10195_ _14360_/D _14427_/Q _14359_/D _06187_/X _14425_/Q VGND VGND VPWR VPWR _14373_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_79_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13954_ _13972_/CLK _13954_/D VGND VGND VPWR VPWR _13954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12905_ _13280_/CLK _12905_/D repeater59/X VGND VGND VPWR VPWR _12905_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13885_ _14210_/CLK _13885_/D VGND VGND VPWR VPWR _13885_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12836_ _14327_/CLK _12836_/D VGND VGND VPWR VPWR hold408/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _13855_/CLK _12767_/D VGND VGND VPWR VPWR hold271/A sky130_fd_sc_hd__dfxtp_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _14615_/CLK _14506_/D VGND VGND VPWR VPWR _14506_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11718_ _11718_/A VGND VGND VPWR VPWR _14051_/D sky130_fd_sc_hd__clkbuf_1
X_12698_ _13283_/CLK _12698_/D VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__dfxtp_1
XFILLER_159_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14437_ _14439_/CLK _14437_/D VGND VGND VPWR VPWR _14437_/Q sky130_fd_sc_hd__dfxtp_1
Xinput11 data_i[19] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_4
X_11649_ _14000_/Q _11516_/X _11653_/S VGND VGND VPWR VPWR _11650_/A sky130_fd_sc_hd__mux2_1
Xinput22 data_i[5] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__buf_4
X_14368_ _14425_/CLK _14368_/D VGND VGND VPWR VPWR _14368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13319_ _14742_/CLK _13319_/D VGND VGND VPWR VPWR _13319_/Q sky130_fd_sc_hd__dfxtp_4
X_14299_ _14705_/CLK _14299_/D VGND VGND VPWR VPWR _14299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08860_ _08860_/A _08860_/B VGND VGND VPWR VPWR _08861_/B sky130_fd_sc_hd__nor2_1
XFILLER_111_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07811_ _07909_/A VGND VGND VPWR VPWR _07811_/X sky130_fd_sc_hd__buf_2
X_08791_ _08791_/A _08791_/B _08791_/C VGND VGND VPWR VPWR _08791_/Y sky130_fd_sc_hd__nand3_1
XFILLER_97_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07742_ _07745_/B VGND VGND VPWR VPWR _07785_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_37_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07673_ _14702_/Q _13115_/Q VGND VGND VPWR VPWR _07675_/C sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_185_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _14733_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09412_ _08556_/B _09411_/Y _09422_/S VGND VGND VPWR VPWR _09413_/A sky130_fd_sc_hd__mux2_1
X_06624_ _12907_/Q _06620_/X _06609_/B VGND VGND VPWR VPWR _06624_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09343_ _13308_/Q _13546_/Q _09343_/S VGND VGND VPWR VPWR _09344_/A sky130_fd_sc_hd__mux2_1
X_06555_ _12890_/Q _06556_/B VGND VGND VPWR VPWR _06557_/A sky130_fd_sc_hd__and2_1
XFILLER_40_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09274_ _09282_/A _09282_/B _07524_/X VGND VGND VPWR VPWR _09274_/X sky130_fd_sc_hd__a21o_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06486_ _12883_/Q _06486_/B VGND VGND VPWR VPWR _06499_/A sky130_fd_sc_hd__nor2_1
X_08225_ _08225_/A _08225_/B VGND VGND VPWR VPWR _08225_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08156_ _08156_/A VGND VGND VPWR VPWR _13357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07107_ _07107_/A _07107_/B _07107_/C VGND VGND VPWR VPWR _07123_/B sky130_fd_sc_hd__or3_1
X_08087_ _12979_/Q _13279_/Q _08095_/S VGND VGND VPWR VPWR _08088_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07038_ _07038_/A _07038_/B VGND VGND VPWR VPWR _07053_/A sky130_fd_sc_hd__and2_1
XFILLER_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08989_ _08989_/A VGND VGND VPWR VPWR _08993_/C sky130_fd_sc_hd__inv_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10951_ _14014_/Q _13980_/Q _13820_/Q _14532_/Q _10921_/X _10922_/X VGND VGND VPWR
+ VPWR _10952_/A sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_176_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _14598_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13670_ _13673_/CLK _13670_/D repeater56/X VGND VGND VPWR VPWR _13670_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10882_ _10882_/A VGND VGND VPWR VPWR _13199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12621_ _12621_/A _12623_/B VGND VGND VPWR VPWR _12621_/X sky130_fd_sc_hd__or2_1
XFILLER_25_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12552_ _11348_/X _14721_/Q _12554_/S VGND VGND VPWR VPWR _12553_/A sky130_fd_sc_hd__mux2_1
X_11503_ _11503_/A VGND VGND VPWR VPWR _13835_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12483_ _12483_/A VGND VGND VPWR VPWR _14672_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_2_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_14222_ _14704_/CLK _14222_/D VGND VGND VPWR VPWR _14222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11434_ _13739_/Q _11438_/B VGND VGND VPWR VPWR _11435_/A sky130_fd_sc_hd__and2_1
X_14153_ _14153_/CLK _14153_/D VGND VGND VPWR VPWR _14153_/Q sky130_fd_sc_hd__dfxtp_1
X_11365_ _12019_/A VGND VGND VPWR VPWR _11365_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_100_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _13945_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13104_ _14530_/CLK hold162/X VGND VGND VPWR VPWR hold467/A sky130_fd_sc_hd__dfxtp_1
XFILLER_113_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10316_ _10312_/A _10309_/Y _10311_/B VGND VGND VPWR VPWR _10317_/B sky130_fd_sc_hd__o21ai_1
X_14084_ _14397_/CLK _14084_/D VGND VGND VPWR VPWR _14084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11296_ _11296_/A VGND VGND VPWR VPWR _13759_/D sky130_fd_sc_hd__clkbuf_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _13294_/CLK _13035_/D VGND VGND VPWR VPWR _13035_/Q sky130_fd_sc_hd__dfxtp_1
X_10247_ _10190_/A _14525_/D _10246_/X VGND VGND VPWR VPWR _10247_/X sky130_fd_sc_hd__a21o_1
XFILLER_67_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10178_ _10178_/A VGND VGND VPWR VPWR _14137_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_167_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _14536_/CLK sky130_fd_sc_hd__clkbuf_16
X_13937_ _13964_/CLK _13937_/D VGND VGND VPWR VPWR _13937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13868_ _14075_/CLK _13868_/D VGND VGND VPWR VPWR _13868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12819_ _13855_/CLK _12819_/D VGND VGND VPWR VPWR hold300/A sky130_fd_sc_hd__dfxtp_1
XFILLER_90_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13799_ _13799_/CLK _13799_/D VGND VGND VPWR VPWR _13799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06340_ _06340_/A VGND VGND VPWR VPWR _14405_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06271_ _13808_/Q _13792_/Q _06273_/S VGND VGND VPWR VPWR _06272_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08010_ _08007_/Y _08008_/X _08003_/A _08004_/Y VGND VGND VPWR VPWR _08010_/X sky130_fd_sc_hd__a211o_1
XFILLER_144_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09961_ _09961_/A VGND VGND VPWR VPWR _12866_/D sky130_fd_sc_hd__clkbuf_1
X_08912_ _08881_/B _08895_/C _08939_/A _08911_/Y VGND VGND VPWR VPWR _08939_/B sky130_fd_sc_hd__o211ai_4
XFILLER_98_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09892_ _13695_/Q _13696_/Q VGND VGND VPWR VPWR _09893_/B sky130_fd_sc_hd__and2_1
XFILLER_98_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08843_ _08944_/A _08843_/B VGND VGND VPWR VPWR _08843_/Y sky130_fd_sc_hd__xnor2_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08774_ _13463_/Q _09563_/B VGND VGND VPWR VPWR _08775_/B sky130_fd_sc_hd__nor2_1
XFILLER_73_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05986_ _14102_/Q _14107_/Q _14108_/Q _14109_/Q VGND VGND VPWR VPWR _05987_/C sky130_fd_sc_hd__or4_1
X_07725_ _07747_/A _07772_/B VGND VGND VPWR VPWR _07726_/B sky130_fd_sc_hd__nand2_1
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_158_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _14327_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_26_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07656_ _07656_/A _07656_/B VGND VGND VPWR VPWR _07657_/B sky130_fd_sc_hd__or2_1
XFILLER_25_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06607_ _12900_/Q _12901_/Q _12902_/Q _06607_/D VGND VGND VPWR VPWR _06620_/B sky130_fd_sc_hd__and4_1
X_07587_ _07583_/B _07583_/C _07583_/A VGND VGND VPWR VPWR _07587_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_159_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09326_ _13300_/Q _13538_/Q _09332_/S VGND VGND VPWR VPWR _09327_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06538_ _06548_/A _06538_/B VGND VGND VPWR VPWR _06538_/Y sky130_fd_sc_hd__xnor2_1
X_09257_ _13549_/Q _09257_/B VGND VGND VPWR VPWR _09264_/A sky130_fd_sc_hd__nand2_1
X_06469_ _06469_/A VGND VGND VPWR VPWR _10339_/A sky130_fd_sc_hd__clkbuf_4
X_08208_ _08208_/A _13427_/Q VGND VGND VPWR VPWR _08250_/C sky130_fd_sc_hd__nor2_1
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09188_ _13538_/Q _09188_/B VGND VGND VPWR VPWR _09188_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08139_ _08135_/B _08137_/Y _08215_/S VGND VGND VPWR VPWR _08140_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11150_ _12645_/B VGND VGND VPWR VPWR _11150_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_161_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10101_ _10179_/S VGND VGND VPWR VPWR _14293_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_89_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11081_ _12585_/A VGND VGND VPWR VPWR _11081_/X sky130_fd_sc_hd__buf_2
XFILLER_150_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10032_ _06082_/X _06256_/X _10032_/S VGND VGND VPWR VPWR _10033_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11983_ _11983_/A VGND VGND VPWR VPWR _14304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_149_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _14714_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13722_ _13722_/CLK hold31/X VGND VGND VPWR VPWR _13722_/Q sky130_fd_sc_hd__dfxtp_1
X_10934_ _12585_/A VGND VGND VPWR VPWR _11208_/A sky130_fd_sc_hd__buf_2
XFILLER_32_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13653_ _13653_/CLK hold61/X VGND VGND VPWR VPWR _14075_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_32_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10865_ _10876_/A VGND VGND VPWR VPWR _10874_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_25_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12604_ _14732_/Q _12616_/A _12604_/C VGND VGND VPWR VPWR _12608_/B sky130_fd_sc_hd__and3_1
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13584_ _14108_/CLK hold166/X VGND VGND VPWR VPWR _13584_/Q sky130_fd_sc_hd__dfxtp_1
X_10796_ _10796_/A VGND VGND VPWR VPWR _13060_/D sky130_fd_sc_hd__clkbuf_1
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12535_ _11313_/X _14713_/Q _12543_/S VGND VGND VPWR VPWR _12536_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12466_ _14664_/Q _12004_/A _12472_/S VGND VGND VPWR VPWR _12467_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14205_ _14209_/CLK _14205_/D VGND VGND VPWR VPWR _14205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11417_ _11417_/A VGND VGND VPWR VPWR _13800_/D sky130_fd_sc_hd__clkbuf_1
X_12397_ _12397_/A VGND VGND VPWR VPWR _14625_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14136_ _14292_/CLK _14136_/D VGND VGND VPWR VPWR hold327/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11348_ _12010_/A VGND VGND VPWR VPWR _11348_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_153_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14067_ _14667_/CLK _14067_/D VGND VGND VPWR VPWR _14067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11279_ _12149_/A _11841_/A VGND VGND VPWR VPWR _12510_/A sky130_fd_sc_hd__or2_4
XFILLER_79_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13018_ _13031_/CLK _13018_/D repeater59/X VGND VGND VPWR VPWR _13018_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_95_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07510_ _07532_/A _07510_/B VGND VGND VPWR VPWR _07510_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08490_ _08490_/A _08490_/B _08489_/X VGND VGND VPWR VPWR _08582_/A sky130_fd_sc_hd__nor3b_1
XFILLER_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07441_ _07442_/A _07443_/A _07442_/B VGND VGND VPWR VPWR _07441_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07372_ _07428_/B _07243_/X _07372_/S VGND VGND VPWR VPWR _07372_/X sky130_fd_sc_hd__mux2_1
X_09111_ _09106_/X _09134_/A _09110_/Y _07307_/X VGND VGND VPWR VPWR _13527_/D sky130_fd_sc_hd__a31o_1
X_06323_ _06323_/A VGND VGND VPWR VPWR _14423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09042_ _09655_/S VGND VGND VPWR VPWR _09051_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06254_ _14393_/D _06254_/B _06254_/C VGND VGND VPWR VPWR _06255_/A sky130_fd_sc_hd__or3_1
XFILLER_117_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold400 hold400/A VGND VGND VPWR VPWR hold400/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06185_ _06185_/A VGND VGND VPWR VPWR _14195_/D sky130_fd_sc_hd__clkbuf_1
Xhold411 hold411/A VGND VGND VPWR VPWR hold411/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold422 hold5/X VGND VGND VPWR VPWR hold422/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold433 hold433/A VGND VGND VPWR VPWR hold433/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold444 hold444/A VGND VGND VPWR VPWR hold444/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold455 hold455/A VGND VGND VPWR VPWR hold455/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold466 hold466/A VGND VGND VPWR VPWR hold466/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold477 hold477/A VGND VGND VPWR VPWR hold477/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold488 hold488/A VGND VGND VPWR VPWR hold488/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09944_ _13496_/Q _13685_/Q _09946_/S VGND VGND VPWR VPWR _09945_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold499 input11/X VGND VGND VPWR VPWR hold499/X sky130_fd_sc_hd__clkbuf_4
XFILLER_58_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _09881_/D _09875_/B VGND VGND VPWR VPWR _13690_/D sky130_fd_sc_hd__nor2_1
XFILLER_97_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08826_ _08826_/A _08826_/B VGND VGND VPWR VPWR _08841_/A sky130_fd_sc_hd__and2_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08757_ _08757_/A _08757_/B VGND VGND VPWR VPWR _08758_/B sky130_fd_sc_hd__and2_1
XFILLER_38_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05969_ _13629_/Q _13638_/Q _13639_/Q _13640_/Q VGND VGND VPWR VPWR _05970_/C sky130_fd_sc_hd__and4_1
XFILLER_57_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _07708_/A _07708_/B VGND VGND VPWR VPWR _07708_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _09563_/B VGND VGND VPWR VPWR _09576_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ _07639_/A VGND VGND VPWR VPWR _13657_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10650_ _10650_/A VGND VGND VPWR VPWR _12678_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09309_ _09309_/A VGND VGND VPWR VPWR _12782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10581_ _13035_/Q _13033_/Q _13030_/Q _06874_/X VGND VGND VPWR VPWR _13030_/D sky130_fd_sc_hd__o31a_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12320_ _14575_/Q _12007_/X _12324_/S VGND VGND VPWR VPWR _12321_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12251_ _11313_/X _14541_/Q _12259_/S VGND VGND VPWR VPWR _12252_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11202_ _14275_/Q _14666_/Q _13773_/Q _14721_/Q _11162_/X _11163_/X VGND VGND VPWR
+ VPWR _11203_/B sky130_fd_sc_hd__mux4_1
XFILLER_119_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12182_ _12182_/A VGND VGND VPWR VPWR _14502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11133_ _11088_/X _11130_/Y _11132_/Y _11095_/X VGND VGND VPWR VPWR _11134_/B sky130_fd_sc_hd__a211o_1
XFILLER_150_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11064_ _13326_/Q _11008_/X _11057_/X _11063_/Y VGND VGND VPWR VPWR _13326_/D sky130_fd_sc_hd__o22a_1
XFILLER_95_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10015_ _10052_/A _13912_/Q VGND VGND VPWR VPWR _10016_/A sky130_fd_sc_hd__xnor2_2
XFILLER_76_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11966_ _14299_/Q _11965_/X _11966_/S VGND VGND VPWR VPWR _11967_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13705_ _14634_/CLK _13705_/D VGND VGND VPWR VPWR hold425/A sky130_fd_sc_hd__dfxtp_2
X_10917_ _11163_/A VGND VGND VPWR VPWR _10918_/A sky130_fd_sc_hd__clkbuf_2
X_14685_ _14687_/CLK hold204/X VGND VGND VPWR VPWR _14685_/Q sky130_fd_sc_hd__dfxtp_1
X_11897_ _11931_/A VGND VGND VPWR VPWR _11948_/S sky130_fd_sc_hd__clkbuf_2
X_13636_ _13653_/CLK hold421/X VGND VGND VPWR VPWR _13636_/Q sky130_fd_sc_hd__dfxtp_1
X_10848_ _13142_/Q _10852_/B VGND VGND VPWR VPWR _10849_/A sky130_fd_sc_hd__and2_1
XFILLER_158_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13567_ _13574_/CLK hold386/X VGND VGND VPWR VPWR _13567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10779_ _13011_/Q _10779_/B VGND VGND VPWR VPWR _10780_/A sky130_fd_sc_hd__and2_1
XFILLER_157_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12518_ _12518_/A VGND VGND VPWR VPWR _14705_/D sky130_fd_sc_hd__clkbuf_1
X_13498_ _13700_/CLK hold433/X VGND VGND VPWR VPWR _13498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12449_ _12449_/A VGND VGND VPWR VPWR _14656_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14119_ _14292_/CLK _14119_/D VGND VGND VPWR VPWR hold253/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07990_ _07995_/A _07990_/B VGND VGND VPWR VPWR _07998_/A sky130_fd_sc_hd__nand2_1
X_06941_ _06932_/A _06932_/B _06935_/A _06934_/X _06950_/A VGND VGND VPWR VPWR _06948_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_68_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09660_ _13711_/Q VGND VGND VPWR VPWR _09767_/A sky130_fd_sc_hd__inv_2
X_06872_ _06861_/X _06869_/X _06870_/Y _06871_/X VGND VGND VPWR VPWR _13013_/D sky130_fd_sc_hd__a31o_1
XFILLER_95_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08611_ _09440_/B _09440_/C _13446_/Q VGND VGND VPWR VPWR _08620_/C sky130_fd_sc_hd__a21oi_1
XFILLER_95_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09591_ _09591_/A VGND VGND VPWR VPWR _12810_/D sky130_fd_sc_hd__clkbuf_2
X_08542_ _08542_/A _08542_/B VGND VGND VPWR VPWR _08542_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08473_ _08545_/S _14245_/Q _08473_/C VGND VGND VPWR VPWR _08473_/X sky130_fd_sc_hd__and3b_1
XFILLER_90_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07424_ _07425_/B _07425_/C _07425_/D _07425_/A VGND VGND VPWR VPWR _07424_/X sky130_fd_sc_hd__a31o_1
XFILLER_149_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07355_ _07355_/A _07367_/B VGND VGND VPWR VPWR _07358_/A sky130_fd_sc_hd__or2_1
XFILLER_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06306_ _06306_/A VGND VGND VPWR VPWR _14187_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07286_ _09099_/A VGND VGND VPWR VPWR _07350_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09025_ _13213_/Q _13442_/Q _09029_/S VGND VGND VPWR VPWR _09026_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06237_ _14089_/Q _12036_/B VGND VGND VPWR VPWR _06238_/A sky130_fd_sc_hd__and2_1
XFILLER_152_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold230 hold230/A VGND VGND VPWR VPWR hold230/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold241 hold241/A VGND VGND VPWR VPWR hold241/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06168_ _06168_/A VGND VGND VPWR VPWR _14171_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold252 hold252/A VGND VGND VPWR VPWR hold252/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold263 hold263/A VGND VGND VPWR VPWR hold263/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold274 hold274/A VGND VGND VPWR VPWR hold274/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold285 hold285/A VGND VGND VPWR VPWR hold285/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_131_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold296 hold296/A VGND VGND VPWR VPWR hold296/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06099_ _13794_/Q _11593_/B VGND VGND VPWR VPWR _06100_/A sky130_fd_sc_hd__and2_1
XFILLER_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09927_ _13488_/Q _13677_/Q _09935_/S VGND VGND VPWR VPWR _09928_/A sky130_fd_sc_hd__mux2_1
X_09858_ _13685_/Q _13686_/Q _09858_/C _09858_/D VGND VGND VPWR VPWR _09873_/C sky130_fd_sc_hd__and4_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08809_ _10306_/A _13511_/D VGND VGND VPWR VPWR _09006_/S sky130_fd_sc_hd__xor2_4
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _09809_/C VGND VGND VPWR VPWR _09836_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _13580_/Q _11828_/B VGND VGND VPWR VPWR _11821_/A sky130_fd_sc_hd__and2_1
XFILLER_65_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11751_/A VGND VGND VPWR VPWR _14066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_80_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _14702_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _10702_/A VGND VGND VPWR VPWR _12929_/D sky130_fd_sc_hd__clkbuf_1
X_14470_ _14539_/CLK _14470_/D VGND VGND VPWR VPWR _14470_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11682_/A VGND VGND VPWR VPWR _14023_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _14333_/CLK hold420/X VGND VGND VPWR VPWR _13421_/Q sky130_fd_sc_hd__dfxtp_1
X_10633_ _14681_/Q _12030_/C _14682_/Q _14688_/Q VGND VGND VPWR VPWR _10634_/A sky130_fd_sc_hd__or4b_1
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13352_ _13353_/CLK _13352_/D VGND VGND VPWR VPWR _13352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10564_ _10564_/A VGND VGND VPWR VPWR _14437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12303_ _12303_/A VGND VGND VPWR VPWR _14567_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13283_ _13283_/CLK _13283_/D repeater59/X VGND VGND VPWR VPWR _13283_/Q sky130_fd_sc_hd__dfrtp_1
X_10495_ _10495_/A _10501_/C VGND VGND VPWR VPWR _10503_/A sky130_fd_sc_hd__nand2_1
X_12234_ _12234_/A VGND VGND VPWR VPWR _14533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12165_ _12165_/A VGND VGND VPWR VPWR _14494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11116_ _12584_/A VGND VGND VPWR VPWR _11116_/X sky130_fd_sc_hd__buf_4
XFILLER_96_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12096_ _12130_/A VGND VGND VPWR VPWR _12147_/S sky130_fd_sc_hd__buf_2
XFILLER_96_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11047_ _11047_/A VGND VGND VPWR VPWR _11047_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 data_i[17] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__buf_6
XFILLER_37_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12998_ _14647_/CLK _12998_/D hold1/X VGND VGND VPWR VPWR _12998_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_91_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14737_ _14737_/CLK _14737_/D VGND VGND VPWR VPWR _14737_/Q sky130_fd_sc_hd__dfxtp_1
X_11949_ _11949_/A VGND VGND VPWR VPWR _14280_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_71_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _13434_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14668_ _14726_/CLK _14668_/D VGND VGND VPWR VPWR _14668_/Q sky130_fd_sc_hd__dfxtp_1
X_13619_ _13619_/CLK _13619_/D repeater57/X VGND VGND VPWR VPWR _13619_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14599_ _14600_/CLK _14599_/D VGND VGND VPWR VPWR _14599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07140_ _07163_/A _07190_/A _07163_/B _07141_/A VGND VGND VPWR VPWR _07142_/A sky130_fd_sc_hd__a22oi_1
XFILLER_158_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07071_ _07072_/A _07072_/B VGND VGND VPWR VPWR _07073_/A sky130_fd_sc_hd__and2_1
XFILLER_146_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06022_ _11819_/A VGND VGND VPWR VPWR _11772_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07973_ _07973_/A _07973_/B VGND VGND VPWR VPWR _07973_/X sky130_fd_sc_hd__or2_1
X_09712_ _09707_/B _09711_/Y _09883_/B VGND VGND VPWR VPWR _09713_/A sky130_fd_sc_hd__mux2_1
X_06924_ _06924_/A _06924_/B _06924_/C _06924_/D VGND VGND VPWR VPWR _06951_/B sky130_fd_sc_hd__or4_1
XFILLER_68_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09643_ _09643_/A VGND VGND VPWR VPWR _12834_/D sky130_fd_sc_hd__clkbuf_1
X_06855_ _13012_/Q _07902_/B VGND VGND VPWR VPWR _06857_/B sky130_fd_sc_hd__xnor2_1
XFILLER_110_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09574_ _09574_/A _09574_/B _09568_/Y _09569_/X VGND VGND VPWR VPWR _09579_/C sky130_fd_sc_hd__or4bb_1
X_06786_ _06786_/A _06786_/B _06786_/C VGND VGND VPWR VPWR _06813_/A sky130_fd_sc_hd__nand3_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _08525_/A VGND VGND VPWR VPWR _08527_/A sky130_fd_sc_hd__clkinv_2
Xclkbuf_leaf_62_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _13525_/CLK sky130_fd_sc_hd__clkbuf_16
X_08456_ _09367_/B _09367_/C _13436_/Q VGND VGND VPWR VPWR _08457_/B sky130_fd_sc_hd__a21oi_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07407_ _13141_/Q _09151_/B _07414_/A _07394_/B VGND VGND VPWR VPWR _07408_/B sky130_fd_sc_hd__o2bb2ai_1
X_08387_ _13090_/Q _13371_/Q _08395_/S VGND VGND VPWR VPWR _08388_/A sky130_fd_sc_hd__mux2_1
X_07338_ _07321_/A _07321_/B _07316_/A _07318_/B _07337_/Y VGND VGND VPWR VPWR _07338_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_149_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07269_ _07267_/S _13655_/Q _07372_/S VGND VGND VPWR VPWR _07269_/X sky130_fd_sc_hd__and3b_1
X_09008_ _13700_/D VGND VGND VPWR VPWR _09655_/S sky130_fd_sc_hd__buf_2
XFILLER_3_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10280_ _10279_/X _10272_/X _10592_/B VGND VGND VPWR VPWR _10281_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13970_ _13972_/CLK _13970_/D VGND VGND VPWR VPWR _13970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12921_ _13039_/CLK _12921_/D VGND VGND VPWR VPWR hold234/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _13727_/CLK _12852_/D VGND VGND VPWR VPWR hold452/A sky130_fd_sc_hd__dfxtp_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _11803_/A VGND VGND VPWR VPWR _14094_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _13574_/CLK _12783_/D VGND VGND VPWR VPWR hold380/A sky130_fd_sc_hd__dfxtp_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _14633_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11734_ _11307_/X _14059_/Q _11736_/S VGND VGND VPWR VPWR _11735_/A sky130_fd_sc_hd__mux2_1
X_14522_ _14555_/CLK _14522_/D VGND VGND VPWR VPWR _14522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14453_ _14610_/CLK _14453_/D VGND VGND VPWR VPWR _14453_/Q sky130_fd_sc_hd__dfxtp_1
X_11665_ _14016_/Q _11459_/X _11667_/S VGND VGND VPWR VPWR _11666_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_4_6_0_clk clkbuf_4_7_0_clk/A VGND VGND VPWR VPWR clkbuf_4_6_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10616_ _10616_/A _10616_/B _10616_/C _10616_/D VGND VGND VPWR VPWR _10616_/X sky130_fd_sc_hd__or4_1
X_13404_ _13606_/CLK hold454/X VGND VGND VPWR VPWR _13404_/Q sky130_fd_sc_hd__dfxtp_1
X_14384_ _14397_/CLK _14384_/D VGND VGND VPWR VPWR hold125/A sky130_fd_sc_hd__dfxtp_1
X_11596_ _13918_/D _13920_/D _11596_/C _13933_/Q VGND VGND VPWR VPWR _11597_/A sky130_fd_sc_hd__or4b_1
X_13335_ _14722_/CLK _13335_/D VGND VGND VPWR VPWR _13335_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10547_ _10547_/A _10547_/B VGND VGND VPWR VPWR _10549_/C sky130_fd_sc_hd__xor2_1
XFILLER_6_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13266_ _13304_/CLK _13266_/D repeater59/X VGND VGND VPWR VPWR _13266_/Q sky130_fd_sc_hd__dfrtp_1
X_10478_ _10468_/X _10471_/B _10469_/A VGND VGND VPWR VPWR _10481_/B sky130_fd_sc_hd__a21oi_1
XFILLER_108_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12217_ _12220_/C _12217_/B VGND VGND VPWR VPWR _14516_/D sky130_fd_sc_hd__nor2_1
XFILLER_142_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13197_ _13617_/CLK _13197_/D VGND VGND VPWR VPWR hold411/A sky130_fd_sc_hd__dfxtp_1
XFILLER_97_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12148_ _12148_/A VGND VGND VPWR VPWR _14488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12079_ _11337_/X _14457_/Q _12085_/S VGND VGND VPWR VPWR _12080_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06640_ _12998_/Q _07802_/A VGND VGND VPWR VPWR _06641_/B sky130_fd_sc_hd__nand2_1
XFILLER_92_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06571_ _06571_/A VGND VGND VPWR VPWR _12891_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_44_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _14435_/CLK sky130_fd_sc_hd__clkbuf_16
X_08310_ _13374_/Q _13375_/Q VGND VGND VPWR VPWR _08317_/D sky130_fd_sc_hd__and2_1
X_09290_ _09285_/A _09286_/X _09289_/Y VGND VGND VPWR VPWR _09290_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_21_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08241_ _08228_/S _08141_/X _08144_/X _08279_/D VGND VGND VPWR VPWR _08243_/B sky130_fd_sc_hd__o211a_1
XANTENNA_14 hold42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_36 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_47 hold473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 input8/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08172_ _08157_/X _08166_/B _08170_/X _08171_/Y VGND VGND VPWR VPWR _13358_/D sky130_fd_sc_hd__a22o_1
XANTENNA_69 _13550_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07123_ _07123_/A _07123_/B _07123_/C VGND VGND VPWR VPWR _07123_/Y sky130_fd_sc_hd__nand3_1
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14754__65 VGND VGND VPWR VPWR _14754__65/HI data_o[28] sky130_fd_sc_hd__conb_1
X_07054_ _07077_/B _07054_/B VGND VGND VPWR VPWR _07055_/B sky130_fd_sc_hd__or2_1
X_06005_ _13577_/Q _13578_/Q _13579_/Q _06005_/D VGND VGND VPWR VPWR _06006_/D sky130_fd_sc_hd__and4_1
XFILLER_88_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07956_ _13273_/Q _07963_/B VGND VGND VPWR VPWR _07957_/B sky130_fd_sc_hd__or2_1
XFILLER_75_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06907_ _07932_/A VGND VGND VPWR VPWR _06907_/X sky130_fd_sc_hd__clkbuf_2
X_07887_ _07859_/A _07859_/B _07859_/C _07859_/D _07886_/Y VGND VGND VPWR VPWR _07887_/Y
+ sky130_fd_sc_hd__o41ai_2
XFILLER_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09626_ _09626_/A VGND VGND VPWR VPWR _12826_/D sky130_fd_sc_hd__clkbuf_1
X_06838_ _06859_/A _07889_/B VGND VGND VPWR VPWR _06838_/X sky130_fd_sc_hd__and2_1
X_09557_ _09559_/B _09557_/B VGND VGND VPWR VPWR _09557_/Y sky130_fd_sc_hd__xnor2_1
X_06769_ _06785_/A _06769_/B VGND VGND VPWR VPWR _06770_/C sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_35_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _12970_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08508_ _08671_/A _08520_/B VGND VGND VPWR VPWR _08509_/B sky130_fd_sc_hd__and2_1
X_09488_ _09510_/A _09509_/A _09484_/A VGND VGND VPWR VPWR _09495_/A sky130_fd_sc_hd__o21a_1
X_08439_ _13435_/Q _09365_/A VGND VGND VPWR VPWR _08440_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11450_ _11523_/S VGND VGND VPWR VPWR _11463_/S sky130_fd_sc_hd__buf_2
XFILLER_7_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10401_ _13520_/Q VGND VGND VPWR VPWR _10429_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_164_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11381_ _11381_/A VGND VGND VPWR VPWR _13784_/D sky130_fd_sc_hd__clkbuf_1
X_13120_ _13657_/CLK _13120_/D VGND VGND VPWR VPWR hold206/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10332_ _13108_/Q _13241_/D _10329_/A VGND VGND VPWR VPWR _10332_/X sky130_fd_sc_hd__a21bo_1
XFILLER_118_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13051_ _13294_/CLK _13051_/D VGND VGND VPWR VPWR hold126/A sky130_fd_sc_hd__dfxtp_1
X_10263_ _10255_/X _14357_/D _10266_/S VGND VGND VPWR VPWR _10263_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12002_ _14310_/Q _12000_/X _12014_/S VGND VGND VPWR VPWR _12003_/A sky130_fd_sc_hd__mux2_1
X_10194_ _10194_/A VGND VGND VPWR VPWR _14360_/D sky130_fd_sc_hd__inv_2
XFILLER_87_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13953_ _13963_/CLK _13953_/D VGND VGND VPWR VPWR _13953_/Q sky130_fd_sc_hd__dfxtp_1
X_12904_ _13280_/CLK _12904_/D hold1/X VGND VGND VPWR VPWR _12904_/Q sky130_fd_sc_hd__dfrtp_1
X_13884_ _14656_/CLK hold502/X VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__dfxtp_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12835_ _14327_/CLK _12835_/D VGND VGND VPWR VPWR hold312/A sky130_fd_sc_hd__dfxtp_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _13565_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _13698_/CLK _12766_/D VGND VGND VPWR VPWR hold262/A sky130_fd_sc_hd__dfxtp_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _14619_/CLK _14505_/D VGND VGND VPWR VPWR _14505_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11717_ _11272_/X _14051_/Q _11725_/S VGND VGND VPWR VPWR _11718_/A sky130_fd_sc_hd__mux2_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12697_ _13027_/CLK _12697_/D VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14436_ _14439_/CLK _14436_/D VGND VGND VPWR VPWR _14436_/Q sky130_fd_sc_hd__dfxtp_1
X_11648_ _11648_/A VGND VGND VPWR VPWR _13999_/D sky130_fd_sc_hd__clkbuf_1
Xinput12 input12/A VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__buf_4
Xinput23 data_i[6] VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__buf_6
XFILLER_128_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14367_ _14425_/CLK _14367_/D VGND VGND VPWR VPWR _14367_/Q sky130_fd_sc_hd__dfxtp_1
X_11579_ _13647_/Q _11585_/B VGND VGND VPWR VPWR _11580_/A sky130_fd_sc_hd__and2_1
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13318_ _14742_/CLK _13318_/D VGND VGND VPWR VPWR _13318_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14298_ _14598_/CLK _14298_/D VGND VGND VPWR VPWR _14298_/Q sky130_fd_sc_hd__dfxtp_1
X_13249_ _14588_/CLK _14588_/Q VGND VGND VPWR VPWR _13249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07810_ _07810_/A VGND VGND VPWR VPWR _13253_/D sky130_fd_sc_hd__clkbuf_1
X_08790_ _08791_/B _08791_/C _08791_/A VGND VGND VPWR VPWR _08790_/X sky130_fd_sc_hd__a21o_1
XFILLER_57_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07741_ _07733_/A _07733_/B _07734_/A VGND VGND VPWR VPWR _07764_/A sky130_fd_sc_hd__a21o_1
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07672_ _13244_/D _13245_/D _07723_/B _13114_/Q VGND VGND VPWR VPWR _07675_/B sky130_fd_sc_hd__and4_1
X_09411_ _09419_/D _09411_/B VGND VGND VPWR VPWR _09411_/Y sky130_fd_sc_hd__xnor2_1
X_06623_ _06623_/A VGND VGND VPWR VPWR _12906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_17_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _14397_/CLK sky130_fd_sc_hd__clkbuf_16
X_09342_ _09342_/A VGND VGND VPWR VPWR _12797_/D sky130_fd_sc_hd__clkbuf_1
X_06554_ _10337_/B _06554_/B _06554_/C VGND VGND VPWR VPWR _06556_/B sky130_fd_sc_hd__and3_1
XFILLER_33_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09273_ _09282_/A _09282_/B VGND VGND VPWR VPWR _09273_/Y sky130_fd_sc_hd__nor2_1
X_06485_ _12883_/Q _06486_/B VGND VGND VPWR VPWR _06493_/B sky130_fd_sc_hd__and2_1
XFILLER_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08224_ _08223_/Y _08214_/B _08211_/A VGND VGND VPWR VPWR _08225_/B sky130_fd_sc_hd__a21oi_1
XFILLER_119_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08155_ _08150_/B _08154_/Y _08215_/S VGND VGND VPWR VPWR _08156_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07106_ _07106_/A _07106_/B VGND VGND VPWR VPWR _07123_/A sky130_fd_sc_hd__nand2_1
XFILLER_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08086_ _08097_/A VGND VGND VPWR VPWR _08095_/S sky130_fd_sc_hd__buf_2
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07037_ _07209_/A VGND VGND VPWR VPWR _07156_/A sky130_fd_sc_hd__buf_2
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08988_ _08988_/A VGND VGND VPWR VPWR _14253_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07939_ _07939_/A _07939_/B _07949_/C VGND VGND VPWR VPWR _07939_/Y sky130_fd_sc_hd__nand3_1
XFILLER_28_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10950_ _14296_/Q _14466_/Q _14222_/Q _14052_/Q _10914_/X _12643_/A VGND VGND VPWR
+ VPWR _10950_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09609_ _13402_/Q _13600_/Q _09609_/S VGND VGND VPWR VPWR _09610_/A sky130_fd_sc_hd__mux2_2
X_10881_ _13157_/Q _10885_/B VGND VGND VPWR VPWR _10882_/A sky130_fd_sc_hd__and2_1
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12620_ _14732_/Q _12616_/B _12619_/X _12617_/X VGND VGND VPWR VPWR _14737_/D sky130_fd_sc_hd__o211a_1
XFILLER_40_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12551_ _12551_/A VGND VGND VPWR VPWR _14720_/D sky130_fd_sc_hd__clkbuf_1
X_11502_ _13835_/Q _11501_/X _11511_/S VGND VGND VPWR VPWR _11503_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12482_ _12484_/A _12484_/B input8/X VGND VGND VPWR VPWR _12483_/A sky130_fd_sc_hd__and3_1
XFILLER_138_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14221_ _14703_/CLK _14221_/D VGND VGND VPWR VPWR _14221_/Q sky130_fd_sc_hd__dfxtp_1
X_11433_ _11433_/A VGND VGND VPWR VPWR _13807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14152_ _14153_/CLK _14152_/D VGND VGND VPWR VPWR _14152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11364_ _11362_/X _11364_/B _11364_/C VGND VGND VPWR VPWR _12019_/A sky130_fd_sc_hd__and3b_4
XFILLER_4_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13103_ _14555_/CLK hold239/X VGND VGND VPWR VPWR hold340/A sky130_fd_sc_hd__dfxtp_1
X_10315_ _10315_/A _10315_/B VGND VGND VPWR VPWR _10317_/A sky130_fd_sc_hd__nand2_1
XFILLER_4_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14083_ _14397_/CLK _14083_/D VGND VGND VPWR VPWR _14083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11295_ _13759_/Q _11294_/X _11295_/S VGND VGND VPWR VPWR _11296_/A sky130_fd_sc_hd__mux2_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ _13039_/CLK _13034_/D VGND VGND VPWR VPWR _13034_/Q sky130_fd_sc_hd__dfxtp_1
X_10246_ _14557_/D _14357_/D VGND VGND VPWR VPWR _10246_/X sky130_fd_sc_hd__and2_1
XFILLER_106_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10177_ _10173_/X _10176_/X _10182_/S VGND VGND VPWR VPWR _10178_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13936_ _14179_/CLK hold86/X VGND VGND VPWR VPWR _13936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13867_ _14075_/CLK _13867_/D VGND VGND VPWR VPWR _13867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12818_ _13855_/CLK _12818_/D VGND VGND VPWR VPWR hold409/A sky130_fd_sc_hd__dfxtp_1
XFILLER_90_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13798_ _13945_/CLK _13798_/D VGND VGND VPWR VPWR _13798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _13702_/CLK _12749_/D VGND VGND VPWR VPWR hold190/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06270_ _06270_/A VGND VGND VPWR VPWR _13953_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14419_ _14732_/CLK _14419_/D VGND VGND VPWR VPWR _14419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09960_ _13503_/Q _13692_/Q _09968_/S VGND VGND VPWR VPWR _09961_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_6_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _14721_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_103_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08911_ _08911_/A _08911_/B _08911_/C VGND VGND VPWR VPWR _08911_/Y sky130_fd_sc_hd__nand3_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _13694_/Q _13695_/Q _09885_/B _13696_/Q VGND VGND VPWR VPWR _09894_/B sky130_fd_sc_hd__a31o_1
XFILLER_97_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _08865_/B _08842_/B VGND VGND VPWR VPWR _08843_/B sky130_fd_sc_hd__or2_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08773_ _13463_/Q _09562_/B VGND VGND VPWR VPWR _08775_/A sky130_fd_sc_hd__and2_1
XFILLER_57_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05985_ _14099_/Q _14100_/Q _14101_/Q _05985_/D VGND VGND VPWR VPWR _05987_/B sky130_fd_sc_hd__or4_1
X_07724_ _07724_/A _07724_/B VGND VGND VPWR VPWR _07726_/A sky130_fd_sc_hd__nor2_1
XFILLER_38_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07655_ _07655_/A _07655_/B VGND VGND VPWR VPWR _07657_/A sky130_fd_sc_hd__nor2_1
XFILLER_81_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06606_ _12901_/Q _06604_/A _06605_/Y VGND VGND VPWR VPWR _12901_/D sky130_fd_sc_hd__a21oi_1
XFILLER_53_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07586_ _13162_/Q _07586_/B VGND VGND VPWR VPWR _07586_/X sky130_fd_sc_hd__or2_1
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09325_ _09325_/A VGND VGND VPWR VPWR _12789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06537_ _06537_/A _06537_/B VGND VGND VPWR VPWR _06538_/B sky130_fd_sc_hd__and2_1
XFILLER_21_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09256_ _09256_/A _09256_/B VGND VGND VPWR VPWR _09261_/C sky130_fd_sc_hd__nand2_1
X_06468_ _06443_/X _06410_/X _06415_/X _06444_/Y VGND VGND VPWR VPWR _06471_/B sky130_fd_sc_hd__o22a_1
X_08207_ _10310_/A _08220_/B _08209_/B VGND VGND VPWR VPWR _08210_/B sky130_fd_sc_hd__and3_1
X_09187_ _09182_/X _09185_/X _09186_/Y _07455_/X VGND VGND VPWR VPWR _13538_/D sky130_fd_sc_hd__a31o_1
X_06399_ _06397_/X _06399_/B VGND VGND VPWR VPWR _06399_/X sky130_fd_sc_hd__and2b_1
XFILLER_135_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08138_ _08303_/A VGND VGND VPWR VPWR _08215_/S sky130_fd_sc_hd__buf_2
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08069_ _12971_/Q _13271_/Q _08073_/S VGND VGND VPWR VPWR _08070_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10100_ _10139_/A _14143_/Q VGND VGND VPWR VPWR _10179_/S sky130_fd_sc_hd__xor2_2
XFILLER_161_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11080_ _14305_/Q _14475_/Q _14231_/Q _14061_/Q _11066_/X _11067_/X VGND VGND VPWR
+ VPWR _11080_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10031_ _10031_/A VGND VGND VPWR VPWR _13969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11982_ _14304_/Q _11981_/X _11982_/S VGND VGND VPWR VPWR _11983_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13721_ _13721_/CLK hold200/X VGND VGND VPWR VPWR _13721_/Q sky130_fd_sc_hd__dfxtp_1
X_10933_ _14745_/Q VGND VGND VPWR VPWR _12585_/A sky130_fd_sc_hd__buf_4
XFILLER_72_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13652_ _14327_/CLK hold401/X VGND VGND VPWR VPWR _13652_/Q sky130_fd_sc_hd__dfxtp_1
X_10864_ _10864_/A VGND VGND VPWR VPWR _13191_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12603_ _12616_/A _12604_/C _12602_/Y VGND VGND VPWR VPWR _14731_/D sky130_fd_sc_hd__a21oi_1
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13583_ _14108_/CLK hold164/X VGND VGND VPWR VPWR _13583_/Q sky130_fd_sc_hd__dfxtp_1
X_10795_ _13018_/Q _10801_/B VGND VGND VPWR VPWR _10796_/A sky130_fd_sc_hd__and2_1
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12534_ _12545_/A VGND VGND VPWR VPWR _12543_/S sky130_fd_sc_hd__buf_2
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12465_ _12465_/A VGND VGND VPWR VPWR _14663_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14204_ _14208_/CLK _14204_/D VGND VGND VPWR VPWR _14204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11416_ _13731_/Q _11416_/B VGND VGND VPWR VPWR _11417_/A sky130_fd_sc_hd__and2_1
X_12396_ hold473/X _12402_/B _12400_/C VGND VGND VPWR VPWR _12397_/A sky130_fd_sc_hd__and3_1
XFILLER_125_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11347_ _13890_/Q _11351_/C _11346_/Y VGND VGND VPWR VPWR _12010_/A sky130_fd_sc_hd__a21oi_4
X_14135_ _14159_/CLK _14135_/D VGND VGND VPWR VPWR hold395/A sky130_fd_sc_hd__dfxtp_1
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14066_ _14615_/CLK _14066_/D VGND VGND VPWR VPWR _14066_/Q sky130_fd_sc_hd__dfxtp_1
X_11278_ _14737_/Q VGND VGND VPWR VPWR _11841_/A sky130_fd_sc_hd__buf_2
XFILLER_140_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10229_ hold497/A _10230_/A _10234_/A VGND VGND VPWR VPWR _14522_/D sky130_fd_sc_hd__a21o_1
X_13017_ _13303_/CLK _13017_/D repeater59/X VGND VGND VPWR VPWR _13017_/Q sky130_fd_sc_hd__dfrtp_1
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__buf_12
XFILLER_94_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13919_ _14042_/CLK _13919_/D VGND VGND VPWR VPWR _13919_/Q sky130_fd_sc_hd__dfxtp_1
X_07440_ _13145_/Q _07444_/A VGND VGND VPWR VPWR _07442_/B sky130_fd_sc_hd__xnor2_2
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07371_ _07326_/X _07365_/X _07369_/X _07370_/Y VGND VGND VPWR VPWR _13139_/D sky130_fd_sc_hd__a22o_1
X_09110_ _09109_/A _09109_/C _09109_/B VGND VGND VPWR VPWR _09110_/Y sky130_fd_sc_hd__o21ai_1
X_06322_ _06321_/X _06216_/A _06322_/S VGND VGND VPWR VPWR _06323_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09041_ _09041_/A VGND VGND VPWR VPWR _12756_/D sky130_fd_sc_hd__clkbuf_1
X_06253_ _14386_/D _14387_/D _14388_/D _14389_/D VGND VGND VPWR VPWR _06254_/C sky130_fd_sc_hd__or4_1
XFILLER_163_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06184_ _14176_/D _06184_/B _06184_/C VGND VGND VPWR VPWR _06185_/A sky130_fd_sc_hd__or3_1
Xhold401 hold401/A VGND VGND VPWR VPWR hold401/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold412 hold412/A VGND VGND VPWR VPWR hold412/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold423 hold423/A VGND VGND VPWR VPWR hold423/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold434 hold434/A VGND VGND VPWR VPWR hold434/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold445 hold445/A VGND VGND VPWR VPWR hold445/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold456 hold456/A VGND VGND VPWR VPWR hold456/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold467 hold467/A VGND VGND VPWR VPWR hold467/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold478 hold8/X VGND VGND VPWR VPWR hold478/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold489 hold489/A VGND VGND VPWR VPWR hold489/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09943_ _09943_/A VGND VGND VPWR VPWR _12858_/D sky130_fd_sc_hd__clkbuf_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _13690_/Q _09872_/A _09855_/X VGND VGND VPWR VPWR _09875_/B sky130_fd_sc_hd__o21ai_1
XFILLER_86_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08825_ _08997_/A VGND VGND VPWR VPWR _08944_/A sky130_fd_sc_hd__buf_2
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05968_ _13641_/Q _13646_/Q _13647_/Q _13648_/Q VGND VGND VPWR VPWR _05970_/B sky130_fd_sc_hd__and4_1
X_08756_ _13459_/Q _13460_/Q _08787_/B VGND VGND VPWR VPWR _08763_/B sky130_fd_sc_hd__o21ai_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07707_ _07733_/A _07705_/Y _07675_/B _07689_/C VGND VGND VPWR VPWR _07710_/B sky130_fd_sc_hd__a211o_1
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08687_ _09555_/B VGND VGND VPWR VPWR _09563_/B sky130_fd_sc_hd__clkbuf_2
X_05899_ hold52/A _13798_/Q _13799_/Q _13802_/Q VGND VGND VPWR VPWR _05904_/C sky130_fd_sc_hd__or4_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ _07616_/Y _07637_/Y _11266_/A VGND VGND VPWR VPWR _07639_/A sky130_fd_sc_hd__mux2_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07569_ _07567_/Y _07568_/X _07526_/X VGND VGND VPWR VPWR _13159_/D sky130_fd_sc_hd__o21bai_1
X_09308_ _13292_/Q _13530_/Q _09310_/S VGND VGND VPWR VPWR _09309_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10580_ _10580_/A VGND VGND VPWR VPWR _13035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09239_ _09241_/B _09239_/B VGND VGND VPWR VPWR _09239_/Y sky130_fd_sc_hd__xnor2_1
X_12250_ _12261_/A VGND VGND VPWR VPWR _12259_/S sky130_fd_sc_hd__buf_2
XFILLER_6_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11201_ _11201_/A VGND VGND VPWR VPWR _11201_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12181_ _14502_/Q _11994_/X _12183_/S VGND VGND VPWR VPWR _12182_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11132_ _11177_/A _11132_/B VGND VGND VPWR VPWR _11132_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11063_ _11108_/A _11063_/B VGND VGND VPWR VPWR _11063_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10014_ _10092_/S VGND VGND VPWR VPWR _14049_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_77_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11965_ _14698_/Q VGND VGND VPWR VPWR _11965_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13704_ _13704_/CLK hold207/X VGND VGND VPWR VPWR _13704_/Q sky130_fd_sc_hd__dfxtp_1
X_10916_ _12584_/A VGND VGND VPWR VPWR _11163_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_45_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14684_ _14688_/CLK hold345/X VGND VGND VPWR VPWR _14684_/Q sky130_fd_sc_hd__dfxtp_1
X_11896_ _12510_/A _12342_/A VGND VGND VPWR VPWR _11931_/A sky130_fd_sc_hd__nor2_8
XFILLER_44_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13635_ _13635_/CLK hold161/X VGND VGND VPWR VPWR _13635_/Q sky130_fd_sc_hd__dfxtp_1
X_10847_ _10847_/A VGND VGND VPWR VPWR _13183_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13566_ _13574_/CLK hold22/X VGND VGND VPWR VPWR _13566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10778_ _10778_/A VGND VGND VPWR VPWR _13052_/D sky130_fd_sc_hd__clkbuf_1
X_12517_ _11288_/X _14705_/Q _12521_/S VGND VGND VPWR VPWR _12518_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13497_ _13700_/CLK hold89/X VGND VGND VPWR VPWR _13497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12448_ _14656_/Q _14513_/Q _12450_/S VGND VGND VPWR VPWR _12449_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12379_ _12379_/A VGND VGND VPWR VPWR _14611_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14118_ _14292_/CLK hold253/X VGND VGND VPWR VPWR _14118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06940_ _06948_/A _06940_/B VGND VGND VPWR VPWR _06950_/A sky130_fd_sc_hd__nor2_1
X_14049_ _14050_/CLK _14049_/D VGND VGND VPWR VPWR _14049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06871_ _06871_/A _07911_/B VGND VGND VPWR VPWR _06871_/X sky130_fd_sc_hd__and2_1
XFILLER_95_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08610_ _13446_/Q _09440_/B _09440_/C VGND VGND VPWR VPWR _08620_/B sky130_fd_sc_hd__and3_1
X_09590_ _13393_/Q _13591_/Q _09598_/S VGND VGND VPWR VPWR _09591_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08541_ _08527_/B _08531_/B _08538_/Y _08525_/A VGND VGND VPWR VPWR _08542_/B sky130_fd_sc_hd__o211a_1
XFILLER_47_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08472_ _08472_/A VGND VGND VPWR VPWR _08545_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_23_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07423_ _13143_/Q _09163_/B VGND VGND VPWR VPWR _07425_/A sky130_fd_sc_hd__xnor2_1
XFILLER_51_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07354_ _13138_/Q _07364_/A _07359_/C VGND VGND VPWR VPWR _07367_/B sky130_fd_sc_hd__and3_1
XFILLER_149_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06305_ _13873_/Q _13857_/Q _10137_/S VGND VGND VPWR VPWR _06306_/A sky130_fd_sc_hd__mux2_1
X_07285_ _07375_/A VGND VGND VPWR VPWR _09099_/A sky130_fd_sc_hd__buf_2
X_09024_ _09024_/A VGND VGND VPWR VPWR _12748_/D sky130_fd_sc_hd__clkbuf_1
X_06236_ _06236_/A VGND VGND VPWR VPWR _14387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold220 hold220/A VGND VGND VPWR VPWR hold220/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06167_ _13857_/Q _11836_/B VGND VGND VPWR VPWR _06168_/A sky130_fd_sc_hd__and2_1
Xhold231 hold231/A VGND VGND VPWR VPWR hold231/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold242 hold242/A VGND VGND VPWR VPWR hold242/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold253 hold253/A VGND VGND VPWR VPWR hold253/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold264 hold264/A VGND VGND VPWR VPWR hold264/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06098_ _06098_/A VGND VGND VPWR VPWR _13939_/D sky130_fd_sc_hd__clkbuf_1
Xhold275 hold275/A VGND VGND VPWR VPWR hold275/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_131_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold286 hold286/A VGND VGND VPWR VPWR hold286/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold297 hold297/A VGND VGND VPWR VPWR hold297/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09926_ _13700_/Q VGND VGND VPWR VPWR _09935_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_58_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _13685_/Q _09851_/X _09856_/Y VGND VGND VPWR VPWR _13685_/D sky130_fd_sc_hd__a21oi_1
XFILLER_100_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ _13473_/D _08808_/B VGND VGND VPWR VPWR _08808_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _09790_/B _09809_/C VGND VGND VPWR VPWR _09791_/B sky130_fd_sc_hd__and2_1
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _08739_/A _08739_/B _08739_/C VGND VGND VPWR VPWR _08739_/X sky130_fd_sc_hd__or3_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11329_/X _14066_/Q _11758_/S VGND VGND VPWR VPWR _11751_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _12886_/Q _10709_/B VGND VGND VPWR VPWR _10702_/A sky130_fd_sc_hd__and2_1
XFILLER_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _14023_/Q _11481_/X _11689_/S VGND VGND VPWR VPWR _11682_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _14696_/CLK hold98/X VGND VGND VPWR VPWR _13420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10632_ _14557_/Q _10630_/X _10631_/X _14556_/Q _14521_/Q VGND VGND VPWR VPWR _14528_/D
+ sky130_fd_sc_hd__a221o_1
X_10563_ _10570_/B _10563_/B VGND VGND VPWR VPWR _10564_/A sky130_fd_sc_hd__and2_1
X_13351_ _13351_/CLK _13351_/D VGND VGND VPWR VPWR _13351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12302_ _14567_/Q _11981_/X _12302_/S VGND VGND VPWR VPWR _12303_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13282_ _13314_/CLK _13282_/D repeater59/X VGND VGND VPWR VPWR _13282_/Q sky130_fd_sc_hd__dfrtp_1
X_10494_ _10495_/A _10501_/C VGND VGND VPWR VPWR _10494_/X sky130_fd_sc_hd__or2_1
XFILLER_5_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12233_ _11288_/X _14533_/Q _12237_/S VGND VGND VPWR VPWR _12234_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12164_ _14494_/Q _11968_/X _12172_/S VGND VGND VPWR VPWR _12165_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11115_ _11186_/A VGND VGND VPWR VPWR _11115_/X sky130_fd_sc_hd__buf_4
X_12095_ _12428_/B _12095_/B VGND VGND VPWR VPWR _12130_/A sky130_fd_sc_hd__nor2_4
XFILLER_122_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11046_ _14603_/Q _14565_/Q _14496_/Q _14448_/Q _11044_/X _11045_/X VGND VGND VPWR
+ VPWR _11047_/A sky130_fd_sc_hd__mux4_1
XFILLER_110_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12997_ _14692_/CLK hold280/X VGND VGND VPWR VPWR hold72/A sky130_fd_sc_hd__dfxtp_1
X_14736_ _14737_/CLK _14736_/D VGND VGND VPWR VPWR _14736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11948_ _14280_/Q _11522_/X _11948_/S VGND VGND VPWR VPWR _11949_/A sky130_fd_sc_hd__mux2_1
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ _14667_/CLK _14667_/D VGND VGND VPWR VPWR _14667_/Q sky130_fd_sc_hd__dfxtp_1
X_11879_ _11879_/A VGND VGND VPWR VPWR _14236_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13618_ _13619_/CLK _13618_/D repeater57/X VGND VGND VPWR VPWR _13618_/Q sky130_fd_sc_hd__dfrtp_1
X_14598_ _14598_/CLK _14598_/D VGND VGND VPWR VPWR _14598_/Q sky130_fd_sc_hd__dfxtp_1
X_13549_ _14555_/CLK _13549_/D _12609_/A VGND VGND VPWR VPWR _13549_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07070_ _07082_/A _07082_/B VGND VGND VPWR VPWR _07072_/B sky130_fd_sc_hd__xnor2_1
X_06021_ _06002_/Y _06006_/X _06020_/X VGND VGND VPWR VPWR _11819_/A sky130_fd_sc_hd__o21ai_4
XFILLER_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07972_ _07972_/A _07972_/B _07972_/C _07970_/C VGND VGND VPWR VPWR _07973_/B sky130_fd_sc_hd__or4b_1
XFILLER_87_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09711_ _09711_/A _09711_/B VGND VGND VPWR VPWR _09711_/Y sky130_fd_sc_hd__xnor2_1
X_06923_ _06932_/A _06923_/B VGND VGND VPWR VPWR _06951_/A sky130_fd_sc_hd__or2_1
XFILLER_101_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09642_ _13417_/Q _13615_/Q _09642_/S VGND VGND VPWR VPWR _09643_/A sky130_fd_sc_hd__mux2_1
X_06854_ _06796_/A _06800_/B _06813_/C _06853_/Y _06769_/B VGND VGND VPWR VPWR _07902_/B
+ sky130_fd_sc_hd__o311a_2
XFILLER_27_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09573_ _13617_/Q _13618_/Q _08787_/B VGND VGND VPWR VPWR _09579_/B sky130_fd_sc_hd__o21ai_1
X_06785_ _06785_/A _06785_/B VGND VGND VPWR VPWR _06786_/C sky130_fd_sc_hd__and2_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _13440_/Q _09401_/B VGND VGND VPWR VPWR _08525_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08455_ _13436_/Q _08490_/A _09367_/C VGND VGND VPWR VPWR _08457_/A sky130_fd_sc_hd__and3_1
XFILLER_51_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07406_ _07414_/B _07414_/C VGND VGND VPWR VPWR _07408_/A sky130_fd_sc_hd__or2_1
XFILLER_23_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08386_ _08397_/A VGND VGND VPWR VPWR _08395_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07337_ _13137_/Q _09118_/B VGND VGND VPWR VPWR _07337_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_109_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07268_ _13171_/Q VGND VGND VPWR VPWR _07372_/S sky130_fd_sc_hd__clkbuf_2
X_06219_ _10208_/S VGND VGND VPWR VPWR _14414_/D sky130_fd_sc_hd__inv_2
X_09007_ _09007_/A VGND VGND VPWR VPWR _14256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07199_ _07184_/X _07198_/Y _07199_/S VGND VGND VPWR VPWR _07200_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09909_ _13480_/Q _13669_/Q _09913_/S VGND VGND VPWR VPWR _09910_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12920_ _13039_/CLK _12920_/D VGND VGND VPWR VPWR hold293/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12851_ _13722_/CLK _12851_/D VGND VGND VPWR VPWR hold83/A sky130_fd_sc_hd__dfxtp_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11802_ _13572_/Q _11806_/B VGND VGND VPWR VPWR _11803_/A sky130_fd_sc_hd__and2_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _13565_/CLK _12782_/D VGND VGND VPWR VPWR hold144/A sky130_fd_sc_hd__dfxtp_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14521_ _14557_/CLK _14521_/D VGND VGND VPWR VPWR _14521_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _11733_/A VGND VGND VPWR VPWR _14058_/D sky130_fd_sc_hd__clkbuf_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _14714_/CLK _14452_/D VGND VGND VPWR VPWR _14452_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _11664_/A VGND VGND VPWR VPWR _14015_/D sky130_fd_sc_hd__clkbuf_1
X_13403_ _13604_/CLK hold342/X VGND VGND VPWR VPWR _13403_/Q sky130_fd_sc_hd__dfxtp_1
X_10615_ _10613_/X _10614_/X _14118_/Q VGND VGND VPWR VPWR _14117_/D sky130_fd_sc_hd__o21a_1
X_14383_ _14413_/CLK _14383_/D VGND VGND VPWR VPWR _14383_/Q sky130_fd_sc_hd__dfxtp_1
X_11595_ _13916_/D _13917_/D _13919_/D _13921_/D VGND VGND VPWR VPWR _11596_/C sky130_fd_sc_hd__or4_1
XFILLER_155_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13334_ _14733_/CLK _13334_/D VGND VGND VPWR VPWR _13334_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_6_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10546_ _12990_/D _10557_/B _10526_/C _10545_/Y VGND VGND VPWR VPWR _10547_/B sky130_fd_sc_hd__a31o_1
XFILLER_10_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13265_ _13265_/CLK _13265_/D repeater59/X VGND VGND VPWR VPWR _13265_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_157_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10477_ _10480_/A _10480_/B VGND VGND VPWR VPWR _10481_/A sky130_fd_sc_hd__xnor2_1
X_12216_ _14123_/Q _12214_/A _12205_/X VGND VGND VPWR VPWR _12217_/B sky130_fd_sc_hd__o21ai_1
X_13196_ _13372_/CLK _13196_/D VGND VGND VPWR VPWR hold457/A sky130_fd_sc_hd__dfxtp_1
XFILLER_96_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12147_ _14488_/Q _12025_/X _12147_/S VGND VGND VPWR VPWR _12148_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12078_ _12078_/A VGND VGND VPWR VPWR _14456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11029_ _14019_/Q _13985_/Q _13825_/Q _14537_/Q _11010_/X _11011_/X VGND VGND VPWR
+ VPWR _11030_/A sky130_fd_sc_hd__mux4_1
XFILLER_92_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06570_ _06565_/B _06569_/Y _06599_/A VGND VGND VPWR VPWR _06571_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14719_ _14720_/CLK _14719_/D VGND VGND VPWR VPWR _14719_/Q sky130_fd_sc_hd__dfxtp_1
X_08240_ _08240_/A VGND VGND VPWR VPWR _13364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_15 hold71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08171_ _08170_/A _08170_/B _07341_/A VGND VGND VPWR VPWR _08171_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_48 hold473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_59 input8/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07122_ _07123_/A _07123_/B _07123_/C VGND VGND VPWR VPWR _07151_/A sky130_fd_sc_hd__a21o_1
XFILLER_158_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07053_ _07053_/A _07053_/B VGND VGND VPWR VPWR _07054_/B sky130_fd_sc_hd__nor2_1
XFILLER_133_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06004_ _13569_/Q _13570_/Q _13571_/Q _13576_/Q VGND VGND VPWR VPWR _06005_/D sky130_fd_sc_hd__and4_1
XFILLER_115_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07955_ _13273_/Q _07955_/B VGND VGND VPWR VPWR _07957_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06906_ _06909_/A _06924_/B VGND VGND VPWR VPWR _06906_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07886_ _07892_/B _07886_/B _07886_/C _07886_/D VGND VGND VPWR VPWR _07886_/Y sky130_fd_sc_hd__nor4_1
XFILLER_28_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09625_ _13409_/Q _13607_/Q _09631_/S VGND VGND VPWR VPWR _09626_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06837_ _06834_/Y _06824_/X _06826_/X _06828_/X _06836_/X VGND VGND VPWR VPWR _06837_/Y
+ sky130_fd_sc_hd__a41oi_1
X_09556_ _09556_/A _09556_/B VGND VGND VPWR VPWR _09557_/B sky130_fd_sc_hd__nand2_1
X_06768_ _06745_/X _06630_/A _06643_/A VGND VGND VPWR VPWR _06769_/B sky130_fd_sc_hd__o21a_1
XFILLER_36_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08507_ _08427_/A _08505_/X _08506_/X _08430_/X _08579_/S _08544_/A VGND VGND VPWR
+ VPWR _08520_/B sky130_fd_sc_hd__mux4_1
X_09487_ _09437_/X _09485_/X _09486_/Y _08764_/X VGND VGND VPWR VPWR _13605_/D sky130_fd_sc_hd__a31o_1
XFILLER_102_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06699_ _06681_/A _06681_/B _06698_/Y VGND VGND VPWR VPWR _06700_/B sky130_fd_sc_hd__o21ai_1
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08438_ _09422_/S VGND VGND VPWR VPWR _09365_/A sky130_fd_sc_hd__buf_2
XFILLER_12_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08369_ _13082_/Q _13363_/Q _08373_/S VGND VGND VPWR VPWR _08370_/A sky130_fd_sc_hd__mux2_1
X_10400_ _10400_/A _10400_/B VGND VGND VPWR VPWR _14216_/D sky130_fd_sc_hd__xnor2_1
X_11380_ _13715_/Q _11382_/B VGND VGND VPWR VPWR _11381_/A sky130_fd_sc_hd__and2_1
XFILLER_164_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10331_ _13109_/Q _13242_/D VGND VGND VPWR VPWR _10334_/A sky130_fd_sc_hd__xor2_1
XFILLER_152_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10262_ _10262_/A VGND VGND VPWR VPWR _14353_/D sky130_fd_sc_hd__clkbuf_1
X_13050_ _13528_/CLK _13050_/D VGND VGND VPWR VPWR hold289/A sky130_fd_sc_hd__dfxtp_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12001_ _12001_/A VGND VGND VPWR VPWR _12014_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_133_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10193_ _10193_/A VGND VGND VPWR VPWR _14359_/D sky130_fd_sc_hd__inv_2
XFILLER_120_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13952_ _13963_/CLK _13952_/D VGND VGND VPWR VPWR _13952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12903_ _13280_/CLK _12903_/D hold1/X VGND VGND VPWR VPWR _12903_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13883_ _14657_/CLK hold60/X VGND VGND VPWR VPWR hold244/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12834_ _14327_/CLK _12834_/D VGND VGND VPWR VPWR hold396/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _13698_/CLK _12765_/D VGND VGND VPWR VPWR hold287/A sky130_fd_sc_hd__dfxtp_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _14615_/CLK _14504_/D VGND VGND VPWR VPWR _14504_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _11766_/S VGND VGND VPWR VPWR _11725_/S sky130_fd_sc_hd__buf_2
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _13304_/CLK _12696_/D VGND VGND VPWR VPWR hold73/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14435_ _14435_/CLK _14435_/D VGND VGND VPWR VPWR _14435_/Q sky130_fd_sc_hd__dfxtp_1
X_11647_ _13999_/Q _11513_/X _11653_/S VGND VGND VPWR VPWR _11648_/A sky130_fd_sc_hd__mux2_1
Xinput13 data_i[20] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__buf_6
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput24 data_i[7] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__buf_8
XFILLER_7_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14366_ _14425_/CLK _14366_/D VGND VGND VPWR VPWR _14366_/Q sky130_fd_sc_hd__dfxtp_1
X_11578_ _11578_/A VGND VGND VPWR VPWR _13870_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13317_ _13565_/CLK hold361/X VGND VGND VPWR VPWR _13317_/Q sky130_fd_sc_hd__dfxtp_1
X_10529_ _10533_/A _10531_/B _10532_/B VGND VGND VPWR VPWR _10537_/A sky130_fd_sc_hd__o21a_1
XFILLER_155_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14297_ _14742_/CLK _14297_/D VGND VGND VPWR VPWR _14297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13248_ _14687_/CLK _14584_/Q VGND VGND VPWR VPWR _13520_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_124_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13179_ _13596_/CLK _13179_/D VGND VGND VPWR VPWR _13212_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07740_ _07740_/A VGND VGND VPWR VPWR _13661_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07671_ _07701_/B _07723_/B _13114_/Q _07701_/A VGND VGND VPWR VPWR _07675_/A sky130_fd_sc_hd__a22oi_2
XFILLER_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09410_ _09419_/C _09403_/B _09409_/Y VGND VGND VPWR VPWR _09411_/B sky130_fd_sc_hd__o21ai_1
XFILLER_53_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06622_ _06620_/X _06622_/B _06622_/C VGND VGND VPWR VPWR _06623_/A sky130_fd_sc_hd__and3b_1
XFILLER_92_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09341_ _13307_/Q _13545_/Q _09343_/S VGND VGND VPWR VPWR _09342_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06553_ _06542_/X _06550_/Y _06552_/Y VGND VGND VPWR VPWR _12889_/D sky130_fd_sc_hd__a21oi_1
XFILLER_40_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09272_ _09272_/A _09272_/B VGND VGND VPWR VPWR _09282_/B sky130_fd_sc_hd__or2_1
X_06484_ _10349_/A _06484_/B _06484_/C VGND VGND VPWR VPWR _06486_/B sky130_fd_sc_hd__and3_1
XFILLER_21_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08223_ _08223_/A VGND VGND VPWR VPWR _08223_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08154_ _08154_/A _08154_/B VGND VGND VPWR VPWR _08154_/Y sky130_fd_sc_hd__xnor2_1
X_07105_ _07105_/A VGND VGND VPWR VPWR _13346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08085_ _08085_/A VGND VGND VPWR VPWR _12702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07036_ _07036_/A VGND VGND VPWR VPWR _13343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08987_ _08972_/X _08986_/Y _08987_/S VGND VGND VPWR VPWR _08988_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_5_0_clk clkbuf_4_5_0_clk/A VGND VGND VPWR VPWR clkbuf_4_5_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07938_ _07939_/A _07939_/B _07949_/C VGND VGND VPWR VPWR _07944_/B sky130_fd_sc_hd__a21o_1
XFILLER_113_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07869_ _06743_/A _06796_/X _07867_/Y _07868_/X VGND VGND VPWR VPWR _13261_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09608_ _09608_/A VGND VGND VPWR VPWR _12818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10880_ _10880_/A VGND VGND VPWR VPWR _13198_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09539_ _09548_/A _09547_/A VGND VGND VPWR VPWR _09539_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12550_ _11343_/X _14720_/Q _12554_/S VGND VGND VPWR VPWR _12551_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11501_ _12004_/A VGND VGND VPWR VPWR _11501_/X sky130_fd_sc_hd__clkbuf_2
X_12481_ _12481_/A VGND VGND VPWR VPWR _14671_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14220_ _14440_/CLK _14220_/D VGND VGND VPWR VPWR _14220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11432_ _13738_/Q _11438_/B VGND VGND VPWR VPWR _11433_/A sky130_fd_sc_hd__and2_1
XFILLER_138_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14151_ _14153_/CLK _14151_/D VGND VGND VPWR VPWR _14151_/Q sky130_fd_sc_hd__dfxtp_1
X_11363_ _13892_/Q _11362_/C _13893_/Q VGND VGND VPWR VPWR _11364_/C sky130_fd_sc_hd__a21o_1
XFILLER_4_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13102_ _14555_/CLK hold250/X VGND VGND VPWR VPWR _13102_/Q sky130_fd_sc_hd__dfxtp_1
X_10314_ _13427_/Q _13514_/D VGND VGND VPWR VPWR _10315_/B sky130_fd_sc_hd__nand2_1
X_14082_ _14082_/CLK _14082_/D VGND VGND VPWR VPWR _14082_/Q sky130_fd_sc_hd__dfxtp_1
X_11294_ _14698_/Q VGND VGND VPWR VPWR _11294_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_152_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ _13294_/CLK _13033_/D VGND VGND VPWR VPWR _13033_/Q sky130_fd_sc_hd__dfxtp_1
X_10245_ _14368_/Q _10230_/X _10237_/A VGND VGND VPWR VPWR _14525_/D sky130_fd_sc_hd__a21o_1
XFILLER_105_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10176_ _10168_/X _14140_/D _10179_/S VGND VGND VPWR VPWR _10176_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13935_ _13972_/CLK _13935_/D VGND VGND VPWR VPWR hold86/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13866_ _14075_/CLK _13866_/D VGND VGND VPWR VPWR _13866_/Q sky130_fd_sc_hd__dfxtp_1
X_12817_ _13855_/CLK _12817_/D VGND VGND VPWR VPWR hold466/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13797_ _13945_/CLK _13797_/D VGND VGND VPWR VPWR _13797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12748_ _13702_/CLK _12748_/D VGND VGND VPWR VPWR hold171/A sky130_fd_sc_hd__dfxtp_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12679_ _14180_/CLK _12679_/D VGND VGND VPWR VPWR _12679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14418_ _14425_/CLK _14418_/D VGND VGND VPWR VPWR _14418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14349_ _14357_/CLK hold472/X VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__dfxtp_1
XFILLER_116_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08910_ _08911_/A _08911_/B _08911_/C VGND VGND VPWR VPWR _08939_/A sky130_fd_sc_hd__a21o_2
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _13695_/Q _09893_/A _09889_/Y VGND VGND VPWR VPWR _13695_/D sky130_fd_sc_hd__a21oi_1
XFILLER_124_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _08841_/A _08841_/B VGND VGND VPWR VPWR _08842_/B sky130_fd_sc_hd__nor2_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _08758_/A _08758_/B _08770_/Y _08771_/X VGND VGND VPWR VPWR _08786_/A sky130_fd_sc_hd__a31oi_2
XFILLER_85_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05984_ _14103_/Q _14104_/Q _14105_/Q _14106_/Q VGND VGND VPWR VPWR _05985_/D sky130_fd_sc_hd__or4_1
XFILLER_84_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07723_ _07723_/A _07723_/B _07723_/C _07745_/B VGND VGND VPWR VPWR _07724_/B sky130_fd_sc_hd__and4_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07654_ _07654_/A _07654_/B VGND VGND VPWR VPWR _07655_/B sky130_fd_sc_hd__nor2_1
XFILLER_41_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06605_ _12901_/Q _06604_/A _06599_/X VGND VGND VPWR VPWR _06605_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07585_ _13162_/Q _09289_/B VGND VGND VPWR VPWR _07585_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09324_ _13299_/Q _13537_/Q _09332_/S VGND VGND VPWR VPWR _09325_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06536_ _06519_/A _06527_/Y _06519_/B _06524_/X _06515_/A VGND VGND VPWR VPWR _06537_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_159_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09255_ _09255_/A _09255_/B VGND VGND VPWR VPWR _09256_/B sky130_fd_sc_hd__and2_1
X_06467_ _06467_/A VGND VGND VPWR VPWR _12881_/D sky130_fd_sc_hd__clkbuf_1
X_08206_ _08206_/A VGND VGND VPWR VPWR _13361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09186_ _09186_/A _09186_/B _09189_/B VGND VGND VPWR VPWR _09186_/Y sky130_fd_sc_hd__nand3_1
X_06398_ _06446_/A _06405_/B _12877_/Q VGND VGND VPWR VPWR _06399_/B sky130_fd_sc_hd__a21o_1
XFILLER_5_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08137_ _08137_/A _08137_/B VGND VGND VPWR VPWR _08137_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_107_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08068_ _08068_/A VGND VGND VPWR VPWR _12694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07019_ _07019_/A _07038_/A VGND VGND VPWR VPWR _07020_/B sky130_fd_sc_hd__or2_1
XFILLER_88_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10030_ _10606_/D _10029_/X _10032_/S VGND VGND VPWR VPWR _10031_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11981_ _14514_/Q VGND VGND VPWR VPWR _11981_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13720_ _13722_/CLK hold36/X VGND VGND VPWR VPWR _13720_/Q sky130_fd_sc_hd__dfxtp_1
X_10932_ _11207_/A VGND VGND VPWR VPWR _10932_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13651_ _14656_/CLK hold328/X VGND VGND VPWR VPWR _13651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10863_ _13149_/Q _10863_/B VGND VGND VPWR VPWR _10864_/A sky130_fd_sc_hd__and2_1
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12602_ _12616_/A _12604_/C _12641_/A VGND VGND VPWR VPWR _12602_/Y sky130_fd_sc_hd__o21ai_1
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13582_ _14275_/CLK hold438/X VGND VGND VPWR VPWR _13582_/Q sky130_fd_sc_hd__dfxtp_1
X_10794_ _10794_/A VGND VGND VPWR VPWR _13059_/D sky130_fd_sc_hd__clkbuf_1
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12533_ _12533_/A VGND VGND VPWR VPWR _14712_/D sky130_fd_sc_hd__clkbuf_1
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12464_ _14663_/Q _14693_/Q _12472_/S VGND VGND VPWR VPWR _12465_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14203_ _14210_/CLK _14203_/D VGND VGND VPWR VPWR _14203_/Q sky130_fd_sc_hd__dfxtp_1
X_11415_ _11415_/A VGND VGND VPWR VPWR _13799_/D sky130_fd_sc_hd__clkbuf_1
X_12395_ _12395_/A VGND VGND VPWR VPWR _14619_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14134_ _14159_/CLK _14134_/D VGND VGND VPWR VPWR hold182/A sky130_fd_sc_hd__dfxtp_1
X_11346_ _13890_/Q _11351_/C _11353_/B VGND VGND VPWR VPWR _11346_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_125_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14065_ _14652_/CLK _14065_/D VGND VGND VPWR VPWR _14065_/Q sky130_fd_sc_hd__dfxtp_1
X_11277_ _14738_/Q VGND VGND VPWR VPWR _12149_/A sky130_fd_sc_hd__buf_2
X_13016_ _13303_/CLK _13016_/D repeater59/X VGND VGND VPWR VPWR _13016_/Q sky130_fd_sc_hd__dfrtp_1
X_10228_ _14521_/D _10236_/B VGND VGND VPWR VPWR _10234_/A sky130_fd_sc_hd__and2_1
XFILLER_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__buf_2
X_10159_ _14294_/D _14140_/D VGND VGND VPWR VPWR _10159_/X sky130_fd_sc_hd__and2_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13918_ _14042_/CLK _13918_/D VGND VGND VPWR VPWR _13918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13849_ _14180_/CLK _13849_/D VGND VGND VPWR VPWR _13849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07370_ _07416_/A _07369_/B _07341_/A VGND VGND VPWR VPWR _07370_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_148_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06321_ _14403_/Q _14395_/Q _06321_/S VGND VGND VPWR VPWR _06321_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06252_ _14390_/D _14391_/D _14392_/D _14413_/D VGND VGND VPWR VPWR _06254_/B sky130_fd_sc_hd__or4_1
X_09040_ _13220_/Q _13449_/Q _09040_/S VGND VGND VPWR VPWR _09041_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06183_ _14169_/D _14170_/D _14171_/D _14172_/D VGND VGND VPWR VPWR _06184_/C sky130_fd_sc_hd__or4_1
Xhold402 hold402/A VGND VGND VPWR VPWR hold402/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold413 hold6/X VGND VGND VPWR VPWR hold413/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold424 hold424/A VGND VGND VPWR VPWR hold424/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold435 hold435/A VGND VGND VPWR VPWR hold435/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold446 hold446/A VGND VGND VPWR VPWR hold446/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold457 hold457/A VGND VGND VPWR VPWR hold457/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_132_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold468 hold7/X VGND VGND VPWR VPWR hold468/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09942_ _13495_/Q _13684_/Q _09946_/S VGND VGND VPWR VPWR _09943_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold479 input12/X VGND VGND VPWR VPWR hold479/X sky130_fd_sc_hd__buf_4
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _13689_/Q _13690_/Q _09873_/C _09873_/D VGND VGND VPWR VPWR _09881_/D sky130_fd_sc_hd__and4_2
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _08824_/A VGND VGND VPWR VPWR _14246_/D sky130_fd_sc_hd__clkbuf_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ _08633_/X _08754_/X _08684_/X VGND VGND VPWR VPWR _13460_/D sky130_fd_sc_hd__a21o_1
X_05967_ _13649_/Q _13650_/Q _13651_/Q _13652_/Q VGND VGND VPWR VPWR _05970_/A sky130_fd_sc_hd__and4_1
XFILLER_85_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07706_ _07675_/B _07689_/C _07733_/A _07705_/Y VGND VGND VPWR VPWR _07733_/B sky130_fd_sc_hd__o211ai_2
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08686_ _09550_/B VGND VGND VPWR VPWR _09555_/B sky130_fd_sc_hd__clkbuf_2
X_05898_ _14622_/Q VGND VGND VPWR VPWR _13119_/D sky130_fd_sc_hd__inv_2
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ _07738_/A _07637_/B VGND VGND VPWR VPWR _07637_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07568_ _07578_/A _07578_/B _07341_/A VGND VGND VPWR VPWR _07568_/X sky130_fd_sc_hd__a21o_1
X_09307_ _09307_/A VGND VGND VPWR VPWR _12781_/D sky130_fd_sc_hd__clkbuf_1
X_06519_ _06519_/A _06519_/B VGND VGND VPWR VPWR _06520_/B sky130_fd_sc_hd__and2_1
XFILLER_70_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07499_ _07499_/A VGND VGND VPWR VPWR _07499_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09238_ _13545_/Q _09289_/B _09234_/A VGND VGND VPWR VPWR _09239_/B sky130_fd_sc_hd__a21oi_1
XFILLER_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09169_ _13536_/Q VGND VGND VPWR VPWR _09177_/A sky130_fd_sc_hd__inv_2
XFILLER_119_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11200_ _14614_/Q _14576_/Q _14507_/Q _14459_/Q _11186_/X _11187_/X VGND VGND VPWR
+ VPWR _11201_/A sky130_fd_sc_hd__mux4_1
XFILLER_134_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12180_ _12180_/A VGND VGND VPWR VPWR _14501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11131_ _14270_/Q _14661_/Q _13768_/Q _14716_/Q _11091_/X _11092_/X VGND VGND VPWR
+ VPWR _11132_/B sky130_fd_sc_hd__mux4_1
XFILLER_150_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11062_ _11017_/X _11059_/Y _11061_/Y _11024_/X VGND VGND VPWR VPWR _11063_/B sky130_fd_sc_hd__a211o_1
XFILLER_89_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10013_ _10052_/A _13911_/Q VGND VGND VPWR VPWR _10092_/S sky130_fd_sc_hd__xor2_2
XFILLER_49_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11964_ _11964_/A VGND VGND VPWR VPWR _14298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13703_ _14251_/CLK _13703_/D VGND VGND VPWR VPWR _13703_/Q sky130_fd_sc_hd__dfxtp_1
X_10915_ _14746_/Q VGND VGND VPWR VPWR _12584_/A sky130_fd_sc_hd__clkbuf_2
X_14683_ _14687_/CLK hold267/X VGND VGND VPWR VPWR _14683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11895_ _11895_/A VGND VGND VPWR VPWR _14244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13634_ _14180_/CLK hold188/X VGND VGND VPWR VPWR _13634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10846_ _13141_/Q _10852_/B VGND VGND VPWR VPWR _10847_/A sky130_fd_sc_hd__and2_1
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13565_ _13565_/CLK hold103/X VGND VGND VPWR VPWR _13565_/Q sky130_fd_sc_hd__dfxtp_1
X_10777_ _13010_/Q _10779_/B VGND VGND VPWR VPWR _10778_/A sky130_fd_sc_hd__and2_1
XFILLER_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12516_ _12516_/A VGND VGND VPWR VPWR _14704_/D sky130_fd_sc_hd__clkbuf_1
X_13496_ _13686_/CLK hold141/X VGND VGND VPWR VPWR _13496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12447_ _12447_/A VGND VGND VPWR VPWR _14655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12378_ _14611_/Q _12000_/X _12386_/S VGND VGND VPWR VPWR _12379_/A sky130_fd_sc_hd__mux2_1
X_14117_ _14292_/CLK _14117_/D VGND VGND VPWR VPWR _14117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11329_ _14693_/Q VGND VGND VPWR VPWR _11329_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14048_ _14210_/CLK _14048_/D VGND VGND VPWR VPWR hold152/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06870_ _06870_/A _06870_/B _06876_/B VGND VGND VPWR VPWR _06870_/Y sky130_fd_sc_hd__nand3_1
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08540_ _08733_/A VGND VGND VPWR VPWR _08542_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08471_ _14249_/Q _14247_/Q _08506_/S VGND VGND VPWR VPWR _08471_/X sky130_fd_sc_hd__mux2_1
X_07422_ _09164_/B VGND VGND VPWR VPWR _09163_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07353_ _13138_/Q _09126_/B VGND VGND VPWR VPWR _07355_/A sky130_fd_sc_hd__nor2_1
XFILLER_148_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06304_ _06304_/A VGND VGND VPWR VPWR _14186_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_137_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07284_ _09086_/B _07284_/B _07283_/X VGND VGND VPWR VPWR _07375_/A sky130_fd_sc_hd__nor3b_1
XFILLER_108_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09023_ _13212_/Q _13441_/Q _09029_/S VGND VGND VPWR VPWR _09024_/A sky130_fd_sc_hd__mux2_1
X_06235_ _14088_/Q _12036_/B VGND VGND VPWR VPWR _06236_/A sky130_fd_sc_hd__and2_1
XFILLER_129_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold210 hold210/A VGND VGND VPWR VPWR hold210/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06166_ _06166_/A VGND VGND VPWR VPWR _14170_/D sky130_fd_sc_hd__clkbuf_1
Xhold221 hold221/A VGND VGND VPWR VPWR hold221/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold232 hold232/A VGND VGND VPWR VPWR hold232/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold243 hold243/A VGND VGND VPWR VPWR hold243/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_117_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold254 hold254/A VGND VGND VPWR VPWR hold254/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06097_ _13793_/Q _11593_/B VGND VGND VPWR VPWR _06098_/A sky130_fd_sc_hd__and2_1
Xhold265 hold265/A VGND VGND VPWR VPWR hold265/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold276 hold276/A VGND VGND VPWR VPWR hold276/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold287 hold287/A VGND VGND VPWR VPWR hold287/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold298 hold298/A VGND VGND VPWR VPWR hold298/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09925_ _09925_/A VGND VGND VPWR VPWR _12850_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ _13685_/Q _09851_/X _09855_/X VGND VGND VPWR VPWR _09856_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_112_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _08807_/A _08826_/A VGND VGND VPWR VPWR _08808_/B sky130_fd_sc_hd__or2_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _09685_/X _09827_/B _09787_/S VGND VGND VPWR VPWR _09790_/B sky130_fd_sc_hd__mux2_1
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06999_ _06999_/A _06999_/B VGND VGND VPWR VPWR _07001_/A sky130_fd_sc_hd__or2_1
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _08739_/A _08739_/B _08739_/C VGND VGND VPWR VPWR _08738_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _08667_/Y _08654_/B _08664_/C _08668_/Y _08662_/B VGND VGND VPWR VPWR _08669_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _13031_/D VGND VGND VPWR VPWR _10709_/B sky130_fd_sc_hd__clkbuf_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11680_ _11691_/A VGND VGND VPWR VPWR _11689_/S sky130_fd_sc_hd__buf_2
XFILLER_53_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10631_ _14527_/Q _14526_/Q VGND VGND VPWR VPWR _10631_/X sky130_fd_sc_hd__or2_1
XFILLER_139_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13350_ _13353_/CLK _13350_/D VGND VGND VPWR VPWR _13350_/Q sky130_fd_sc_hd__dfxtp_1
X_10562_ _10562_/A _10562_/B _10562_/C VGND VGND VPWR VPWR _10563_/B sky130_fd_sc_hd__or3_1
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12301_ _12301_/A VGND VGND VPWR VPWR _14566_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13281_ _13314_/CLK _13281_/D repeater59/X VGND VGND VPWR VPWR _13281_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10493_ _10493_/A _10488_/B VGND VGND VPWR VPWR _10498_/A sky130_fd_sc_hd__or2b_1
XFILLER_154_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12232_ _12232_/A VGND VGND VPWR VPWR _14532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12163_ _12185_/A VGND VGND VPWR VPWR _12172_/S sky130_fd_sc_hd__buf_2
XFILLER_107_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11114_ _11185_/A VGND VGND VPWR VPWR _11179_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_96_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12094_ _12094_/A VGND VGND VPWR VPWR _14464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11045_ _11153_/A VGND VGND VPWR VPWR _11045_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12996_ _13296_/CLK hold49/X VGND VGND VPWR VPWR hold500/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14735_ _14746_/CLK _14735_/D VGND VGND VPWR VPWR _14735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11947_ _11947_/A VGND VGND VPWR VPWR _14279_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14666_ _14667_/CLK _14666_/D VGND VGND VPWR VPWR _14666_/Q sky130_fd_sc_hd__dfxtp_1
X_11878_ _14236_/Q _11497_/X _11886_/S VGND VGND VPWR VPWR _11879_/A sky130_fd_sc_hd__mux2_1
X_13617_ _13617_/CLK _13617_/D repeater57/X VGND VGND VPWR VPWR _13617_/Q sky130_fd_sc_hd__dfrtp_1
X_10829_ _13134_/Q _10893_/A VGND VGND VPWR VPWR _10830_/A sky130_fd_sc_hd__and2_1
X_14597_ _14749_/CLK _14597_/D VGND VGND VPWR VPWR _14597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13548_ _14082_/CLK _13548_/D _12609_/A VGND VGND VPWR VPWR _13548_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13479_ _14251_/CLK hold116/X VGND VGND VPWR VPWR _13479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06020_ _06007_/X _06008_/X _06012_/X _06019_/Y VGND VGND VPWR VPWR _06020_/X sky130_fd_sc_hd__a31o_1
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07971_ _06793_/A _07969_/Y _07970_/X _07940_/X VGND VGND VPWR VPWR _13275_/D sky130_fd_sc_hd__a31o_1
XFILLER_114_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09710_ _09697_/A _09696_/A _09709_/X VGND VGND VPWR VPWR _09711_/B sky130_fd_sc_hd__a21o_1
XFILLER_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06922_ _13018_/Q _06954_/A VGND VGND VPWR VPWR _06923_/B sky130_fd_sc_hd__nor2_1
XFILLER_113_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09641_ _09641_/A VGND VGND VPWR VPWR _12833_/D sky130_fd_sc_hd__clkbuf_1
X_06853_ _06747_/Y _06852_/Y _06745_/X VGND VGND VPWR VPWR _06853_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09572_ _09502_/X _09570_/Y _09571_/X _09506_/X VGND VGND VPWR VPWR _13618_/D sky130_fd_sc_hd__a31o_1
X_06784_ _06863_/A _06783_/X _06769_/B VGND VGND VPWR VPWR _06785_/B sky130_fd_sc_hd__o21a_1
X_08523_ _08523_/A VGND VGND VPWR VPWR _09401_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_24_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08454_ _09367_/B _09367_/C VGND VGND VPWR VPWR _08454_/X sky130_fd_sc_hd__and2_1
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07405_ _09153_/B _09153_/C _13142_/Q VGND VGND VPWR VPWR _07414_/C sky130_fd_sc_hd__a21oi_1
XFILLER_11_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08385_ _08385_/A VGND VGND VPWR VPWR _12725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07336_ _09118_/B VGND VGND VPWR VPWR _07356_/B sky130_fd_sc_hd__clkbuf_2
X_07267_ _13659_/Q _13657_/Q _07267_/S VGND VGND VPWR VPWR _07267_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09006_ _09003_/Y _13473_/D _09006_/S VGND VGND VPWR VPWR _09007_/A sky130_fd_sc_hd__mux2_1
X_06218_ _06322_/S VGND VGND VPWR VPWR _10208_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_152_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07198_ _07209_/A _07198_/B VGND VGND VPWR VPWR _07198_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_117_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06149_ _10121_/S VGND VGND VPWR VPWR _14197_/D sky130_fd_sc_hd__inv_2
XFILLER_78_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09908_ _09908_/A VGND VGND VPWR VPWR _12842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09839_ _09839_/A _09839_/B VGND VGND VPWR VPWR _09842_/A sky130_fd_sc_hd__nor2_1
XFILLER_58_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12850_ _13721_/CLK _12850_/D VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11801_ _11801_/A VGND VGND VPWR VPWR _14093_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _13574_/CLK _12781_/D VGND VGND VPWR VPWR hold192/A sky130_fd_sc_hd__dfxtp_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14520_ _14530_/CLK hold120/X VGND VGND VPWR VPWR _14520_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _11304_/X _14058_/Q _11736_/S VGND VGND VPWR VPWR _11733_/A sky130_fd_sc_hd__mux2_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14602_/CLK _14451_/D VGND VGND VPWR VPWR _14451_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _14015_/Q _11456_/X _11667_/S VGND VGND VPWR VPWR _11664_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _13621_/CLK hold463/X VGND VGND VPWR VPWR _13402_/Q sky130_fd_sc_hd__dfxtp_1
X_10614_ _14289_/Q _14146_/Q _14154_/Q hold429/A VGND VGND VPWR VPWR _10614_/X sky130_fd_sc_hd__or4_1
X_14382_ _14397_/CLK hold230/X VGND VGND VPWR VPWR _14382_/Q sky130_fd_sc_hd__dfxtp_1
X_11594_ _11594_/A VGND VGND VPWR VPWR _13934_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13333_ _14733_/CLK _13333_/D VGND VGND VPWR VPWR _13333_/Q sky130_fd_sc_hd__dfxtp_4
X_10545_ _10545_/A VGND VGND VPWR VPWR _10545_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_130_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _14042_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13264_ _13264_/CLK _13264_/D repeater59/X VGND VGND VPWR VPWR _13264_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_155_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10476_ _10476_/A _10476_/B VGND VGND VPWR VPWR _10480_/B sky130_fd_sc_hd__xor2_1
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12215_ _14122_/Q _14123_/Q _12215_/C VGND VGND VPWR VPWR _12220_/C sky130_fd_sc_hd__and3_1
XFILLER_124_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13195_ _13606_/CLK _13195_/D VGND VGND VPWR VPWR hold514/A sky130_fd_sc_hd__dfxtp_1
X_12146_ _12146_/A VGND VGND VPWR VPWR _14487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12077_ _11329_/X _14456_/Q _12085_/S VGND VGND VPWR VPWR _12078_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11028_ _14301_/Q _14471_/Q _14227_/Q _14057_/Q _10993_/X _10995_/X VGND VGND VPWR
+ VPWR _11028_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12979_ _13280_/CLK hold285/X VGND VGND VPWR VPWR _12979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14718_ _14720_/CLK _14718_/D VGND VGND VPWR VPWR _14718_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14649_ _14703_/CLK _14649_/D VGND VGND VPWR VPWR _14649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_16 hold42/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_27 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_38 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08170_ _08170_/A _08170_/B VGND VGND VPWR VPWR _08170_/X sky130_fd_sc_hd__or2_1
XANTENNA_49 _14729_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07121_ _07121_/A _07121_/B VGND VGND VPWR VPWR _07123_/C sky130_fd_sc_hd__xnor2_1
XFILLER_146_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_121_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _13855_/CLK sky130_fd_sc_hd__clkbuf_16
X_07052_ _07053_/A _07053_/B VGND VGND VPWR VPWR _07077_/B sky130_fd_sc_hd__and2_1
XFILLER_115_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06003_ _13565_/Q _13566_/Q _13567_/Q _13568_/Q VGND VGND VPWR VPWR _06006_/C sky130_fd_sc_hd__and4_1
XFILLER_126_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07954_ _07909_/X _07952_/X _07953_/Y _07940_/X VGND VGND VPWR VPWR _13272_/D sky130_fd_sc_hd__a31o_1
XFILLER_29_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06905_ _06909_/A _06924_/B VGND VGND VPWR VPWR _06905_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_188_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _14725_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07885_ _07885_/A _07885_/B _07885_/C _07885_/D VGND VGND VPWR VPWR _07886_/B sky130_fd_sc_hd__or4_1
XFILLER_110_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09624_ _09624_/A VGND VGND VPWR VPWR _12825_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06836_ _06895_/A VGND VGND VPWR VPWR _06836_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09555_ _13616_/Q _09555_/B VGND VGND VPWR VPWR _09559_/B sky130_fd_sc_hd__xnor2_1
XFILLER_71_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06767_ _06782_/A _06767_/B VGND VGND VPWR VPWR _06785_/A sky130_fd_sc_hd__or2_1
XFILLER_36_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08506_ _14251_/Q _14249_/Q _08506_/S VGND VGND VPWR VPWR _08506_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09486_ _09510_/A _09509_/A VGND VGND VPWR VPWR _09486_/Y sky130_fd_sc_hd__nand2_1
X_06698_ _13000_/Q _07821_/B VGND VGND VPWR VPWR _06698_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08437_ _13469_/Q VGND VGND VPWR VPWR _09422_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08368_ _08368_/A VGND VGND VPWR VPWR _12717_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07319_ _13135_/Q _09113_/B VGND VGND VPWR VPWR _07320_/A sky130_fd_sc_hd__and2_1
X_08299_ _13372_/Q _08294_/X _08298_/X VGND VGND VPWR VPWR _08299_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_112_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _13372_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10330_ _13749_/Q _10330_/B VGND VGND VPWR VPWR _13242_/D sky130_fd_sc_hd__xnor2_4
XFILLER_164_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10261_ _10256_/X _10260_/X _14555_/D VGND VGND VPWR VPWR _10262_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12000_ _14693_/Q VGND VGND VPWR VPWR _12000_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10192_ _10230_/A VGND VGND VPWR VPWR _14521_/D sky130_fd_sc_hd__inv_2
XFILLER_87_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_179_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _14705_/CLK sky130_fd_sc_hd__clkbuf_16
X_13951_ _13963_/CLK _13951_/D VGND VGND VPWR VPWR _13951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12902_ _13274_/CLK _12902_/D hold1/X VGND VGND VPWR VPWR _12902_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13882_ _14657_/CLK hold244/X VGND VGND VPWR VPWR hold236/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12833_ _14327_/CLK _12833_/D VGND VGND VPWR VPWR hold357/A sky130_fd_sc_hd__dfxtp_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _13700_/CLK _12764_/D VGND VGND VPWR VPWR hold277/A sky130_fd_sc_hd__dfxtp_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14503_ _14610_/CLK _14503_/D VGND VGND VPWR VPWR _14503_/Q sky130_fd_sc_hd__dfxtp_1
X_11715_ _11749_/A VGND VGND VPWR VPWR _11766_/S sky130_fd_sc_hd__buf_2
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _13304_/CLK _12695_/D VGND VGND VPWR VPWR hold189/A sky130_fd_sc_hd__dfxtp_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14434_ _14439_/CLK _14434_/D VGND VGND VPWR VPWR _14434_/Q sky130_fd_sc_hd__dfxtp_1
X_11646_ _11646_/A VGND VGND VPWR VPWR _13998_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput14 data_i[21] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_2
Xinput25 data_i[8] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14365_ _14425_/CLK _14365_/D VGND VGND VPWR VPWR hold497/A sky130_fd_sc_hd__dfxtp_1
X_11577_ _13646_/Q _11585_/B VGND VGND VPWR VPWR _11578_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_103_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _13700_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_156_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13316_ _14098_/CLK hold332/X VGND VGND VPWR VPWR _13316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10528_ _14430_/D _10557_/B _10526_/C VGND VGND VPWR VPWR _10532_/B sky130_fd_sc_hd__a21o_1
XFILLER_156_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14296_ _14703_/CLK _14296_/D VGND VGND VPWR VPWR _14296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13247_ _14687_/CLK _13247_/D VGND VGND VPWR VPWR _13519_/D sky130_fd_sc_hd__dfxtp_1
X_10459_ _10460_/A _10456_/X _10476_/A VGND VGND VPWR VPWR _10463_/A sky130_fd_sc_hd__o21ba_1
XFILLER_124_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13178_ _13596_/CLK _13178_/D VGND VGND VPWR VPWR hold437/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12129_ _12129_/A VGND VGND VPWR VPWR _14479_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07670_ _07688_/A _07688_/B VGND VGND VPWR VPWR _07689_/A sky130_fd_sc_hd__xnor2_1
XFILLER_37_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06621_ _12905_/Q _06616_/A _12906_/Q VGND VGND VPWR VPWR _06622_/C sky130_fd_sc_hd__a21o_1
XFILLER_80_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09340_ _09340_/A VGND VGND VPWR VPWR _12796_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06552_ _06609_/B _06552_/B VGND VGND VPWR VPWR _06552_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09271_ _13551_/Q _09271_/B VGND VGND VPWR VPWR _09272_/B sky130_fd_sc_hd__nor2_1
X_06483_ _06543_/A _10339_/A _12671_/Q _06502_/A VGND VGND VPWR VPWR _06484_/C sky130_fd_sc_hd__a31o_1
X_08222_ _08222_/A _08234_/A VGND VGND VPWR VPWR _08225_/A sky130_fd_sc_hd__or2_1
X_08153_ _08137_/A _08136_/A _08152_/X VGND VGND VPWR VPWR _08154_/B sky130_fd_sc_hd__a21o_1
XFILLER_119_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07104_ _07079_/Y _07102_/Y _07199_/S VGND VGND VPWR VPWR _07105_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08084_ _12978_/Q _13278_/Q _08084_/S VGND VGND VPWR VPWR _08085_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07035_ _07020_/Y _07034_/Y _10647_/A VGND VGND VPWR VPWR _07036_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08986_ _08997_/A _08986_/B VGND VGND VPWR VPWR _08986_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07937_ _07944_/A _07937_/B VGND VGND VPWR VPWR _07949_/C sky130_fd_sc_hd__nand2_1
XFILLER_29_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07868_ _07885_/C _07892_/A _07866_/X _06976_/A VGND VGND VPWR VPWR _07868_/X sky130_fd_sc_hd__o31a_1
XFILLER_84_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09607_ _13401_/Q _13599_/Q _09609_/S VGND VGND VPWR VPWR _09608_/A sky130_fd_sc_hd__mux2_2
X_06819_ _06820_/A _06820_/B _06820_/C VGND VGND VPWR VPWR _06819_/X sky130_fd_sc_hd__a21o_1
XFILLER_73_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07799_ _07799_/A VGND VGND VPWR VPWR _13665_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09538_ _13613_/Q _09542_/B VGND VGND VPWR VPWR _09547_/A sky130_fd_sc_hd__xor2_1
XFILLER_24_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09469_ _09477_/A _09468_/B _08542_/A VGND VGND VPWR VPWR _09469_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11500_ _11500_/A VGND VGND VPWR VPWR _13834_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12480_ _14671_/Q _12025_/A _12480_/S VGND VGND VPWR VPWR _12481_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11431_ _11431_/A VGND VGND VPWR VPWR _13806_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14150_ _14153_/CLK _14150_/D VGND VGND VPWR VPWR _14150_/Q sky130_fd_sc_hd__dfxtp_1
X_11362_ _13892_/Q _13893_/Q _11362_/C VGND VGND VPWR VPWR _11362_/X sky130_fd_sc_hd__and3_1
XFILLER_153_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13101_ _14555_/CLK hold446/X VGND VGND VPWR VPWR hold469/A sky130_fd_sc_hd__dfxtp_1
XFILLER_153_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10313_ _13427_/Q _13514_/D VGND VGND VPWR VPWR _10315_/A sky130_fd_sc_hd__or2_1
XFILLER_4_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14081_ _14397_/CLK _14081_/D VGND VGND VPWR VPWR _14081_/Q sky130_fd_sc_hd__dfxtp_1
X_11293_ _11293_/A VGND VGND VPWR VPWR _13758_/D sky130_fd_sc_hd__clkbuf_1
X_13032_ _13294_/CLK hold506/X VGND VGND VPWR VPWR _13032_/Q sky130_fd_sc_hd__dfxtp_1
X_10244_ _10244_/A VGND VGND VPWR VPWR _14527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10175_ _10175_/A VGND VGND VPWR VPWR _14136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13934_ _13964_/CLK _13934_/D VGND VGND VPWR VPWR _13934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13865_ _14075_/CLK _13865_/D VGND VGND VPWR VPWR _13865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12816_ _13653_/CLK _12816_/D VGND VGND VPWR VPWR hold142/A sky130_fd_sc_hd__dfxtp_1
XFILLER_90_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13796_ _13945_/CLK _13796_/D VGND VGND VPWR VPWR _13796_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _13702_/CLK _12747_/D VGND VGND VPWR VPWR hold195/A sky130_fd_sc_hd__dfxtp_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ _14413_/CLK _12678_/D VGND VGND VPWR VPWR _12678_/Q sky130_fd_sc_hd__dfxtp_1
X_11629_ _11629_/A VGND VGND VPWR VPWR _13990_/D sky130_fd_sc_hd__clkbuf_1
X_14417_ _14732_/CLK _14417_/D VGND VGND VPWR VPWR _14417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14348_ _14357_/CLK hold439/X VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__dfxtp_1
XFILLER_144_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14279_ _14725_/CLK _14279_/D VGND VGND VPWR VPWR _14279_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _08841_/A _08841_/B VGND VGND VPWR VPWR _08865_/B sky130_fd_sc_hd__and2_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _13459_/Q _13460_/Q _13461_/Q _13462_/Q _09563_/B VGND VGND VPWR VPWR _08771_/X
+ sky130_fd_sc_hd__o41a_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05983_ hold77/A _14094_/Q _05983_/C VGND VGND VPWR VPWR _05987_/A sky130_fd_sc_hd__or3_1
XFILLER_111_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07722_ _07745_/A _07772_/A _07745_/B _07723_/A VGND VGND VPWR VPWR _07724_/A sky130_fd_sc_hd__a22oi_1
X_07653_ _07654_/A _07654_/B VGND VGND VPWR VPWR _07655_/A sky130_fd_sc_hd__and2_1
XFILLER_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06604_ _06604_/A _06604_/B VGND VGND VPWR VPWR _12900_/D sky130_fd_sc_hd__nor2_1
XFILLER_92_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07584_ _07570_/X _07582_/X _07583_/Y _07575_/X VGND VGND VPWR VPWR _13161_/D sky130_fd_sc_hd__a31o_1
XFILLER_41_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09323_ _09323_/A VGND VGND VPWR VPWR _09332_/S sky130_fd_sc_hd__clkbuf_2
X_06535_ _06535_/A _06535_/B VGND VGND VPWR VPWR _06548_/A sky130_fd_sc_hd__or2_1
XFILLER_40_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09254_ _13547_/Q _13548_/Q _09284_/B VGND VGND VPWR VPWR _09261_/B sky130_fd_sc_hd__o21ai_1
X_06466_ _06462_/B _06465_/Y _06622_/B VGND VGND VPWR VPWR _06467_/A sky130_fd_sc_hd__mux2_1
X_08205_ _08201_/B _08204_/Y _08215_/S VGND VGND VPWR VPWR _08206_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09185_ _09186_/A _09186_/B _09189_/B VGND VGND VPWR VPWR _09185_/X sky130_fd_sc_hd__a21o_1
X_06397_ _06446_/A _12877_/Q _06405_/B VGND VGND VPWR VPWR _06397_/X sky130_fd_sc_hd__and3_1
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08136_ _08136_/A _08136_/B VGND VGND VPWR VPWR _08137_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08067_ _12970_/Q _13270_/Q _08073_/S VGND VGND VPWR VPWR _08068_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07018_ _07040_/A _07031_/A _07045_/C VGND VGND VPWR VPWR _07038_/A sky130_fd_sc_hd__and3_1
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08969_ _08970_/A _08970_/B _08970_/C VGND VGND VPWR VPWR _08971_/A sky130_fd_sc_hd__a21oi_1
XFILLER_124_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11980_ _11980_/A VGND VGND VPWR VPWR _14303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10931_ _12590_/A VGND VGND VPWR VPWR _11207_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13650_ _14327_/CLK hold408/X VGND VGND VPWR VPWR _13650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10862_ _10862_/A VGND VGND VPWR VPWR _13190_/D sky130_fd_sc_hd__clkbuf_1
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12601_ _14731_/Q VGND VGND VPWR VPWR _12616_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13581_ _14275_/CLK hold375/X VGND VGND VPWR VPWR _13581_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10793_ _13017_/Q _10801_/B VGND VGND VPWR VPWR _10794_/A sky130_fd_sc_hd__and2_1
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12532_ _11310_/X _14712_/Q _12532_/S VGND VGND VPWR VPWR _12533_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12463_ _12463_/A VGND VGND VPWR VPWR _12472_/S sky130_fd_sc_hd__buf_2
X_14202_ _14210_/CLK _14202_/D VGND VGND VPWR VPWR _14202_/Q sky130_fd_sc_hd__dfxtp_1
X_11414_ _13730_/Q _11416_/B VGND VGND VPWR VPWR _11415_/A sky130_fd_sc_hd__and2_1
X_12394_ _14619_/Q _12025_/X _12394_/S VGND VGND VPWR VPWR _12395_/A sky130_fd_sc_hd__mux2_1
X_14133_ _14292_/CLK hold393/X VGND VGND VPWR VPWR hold243/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11345_ _11345_/A VGND VGND VPWR VPWR _13772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14064_ _14652_/CLK _14064_/D VGND VGND VPWR VPWR _14064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11276_ _11712_/B _12582_/A _14736_/Q VGND VGND VPWR VPWR _12150_/A sky130_fd_sc_hd__or3b_4
XFILLER_98_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13015_ _13303_/CLK _13015_/D repeater59/X VGND VGND VPWR VPWR _13015_/Q sky130_fd_sc_hd__dfrtp_1
X_10227_ _10236_/B VGND VGND VPWR VPWR _14357_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10158_ _14151_/Q _10143_/X _10150_/A VGND VGND VPWR VPWR _14286_/D sky130_fd_sc_hd__a21o_1
XFILLER_95_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3 rst_n VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10089_ _10081_/X _13908_/D _10092_/S VGND VGND VPWR VPWR _10089_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13917_ _14042_/CLK _13917_/D VGND VGND VPWR VPWR _13917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13848_ _14180_/CLK _13848_/D VGND VGND VPWR VPWR _13848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13779_ _14633_/CLK _13779_/D VGND VGND VPWR VPWR hold203/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06320_ _14186_/D _14187_/D _06316_/X _06319_/Y VGND VGND VPWR VPWR _14193_/D sky130_fd_sc_hd__a31o_1
XFILLER_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06251_ _06249_/X _06250_/X _12036_/B VGND VGND VPWR VPWR _14413_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_4_4_0_clk clkbuf_4_5_0_clk/A VGND VGND VPWR VPWR clkbuf_4_4_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06182_ _14173_/D _14174_/D _14175_/D _14196_/D VGND VGND VPWR VPWR _06184_/B sky130_fd_sc_hd__or4_1
XFILLER_129_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold403 hold44/X VGND VGND VPWR VPWR hold403/X sky130_fd_sc_hd__clkbuf_1
Xhold414 hold414/A VGND VGND VPWR VPWR hold414/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_128_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold425 hold425/A VGND VGND VPWR VPWR hold425/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold436 hold436/A VGND VGND VPWR VPWR hold436/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_143_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold447 hold447/A VGND VGND VPWR VPWR hold447/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold458 hold458/A VGND VGND VPWR VPWR hold458/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_143_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold469 hold469/A VGND VGND VPWR VPWR hold469/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09941_ _09941_/A VGND VGND VPWR VPWR _12857_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _09872_/A _09872_/B VGND VGND VPWR VPWR _13689_/D sky130_fd_sc_hd__nor2_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08823_ _08808_/Y _08822_/Y _11268_/A VGND VGND VPWR VPWR _08824_/A sky130_fd_sc_hd__mux2_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08754_ _08757_/B _08754_/B VGND VGND VPWR VPWR _08754_/X sky130_fd_sc_hd__xor2_1
X_05966_ _14075_/D _13622_/Q _13623_/Q _13624_/Q VGND VGND VPWR VPWR _05966_/X sky130_fd_sc_hd__and4_1
XFILLER_85_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07705_ _07705_/A _07705_/B _07705_/C VGND VGND VPWR VPWR _07705_/Y sky130_fd_sc_hd__nand3_1
XFILLER_26_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08685_ _08633_/X _08675_/Y _08684_/X VGND VGND VPWR VPWR _13451_/D sky130_fd_sc_hd__a21o_1
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05897_ _13747_/Q VGND VGND VPWR VPWR _13240_/D sky130_fd_sc_hd__clkinv_2
XFILLER_93_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_92_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _14250_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _07659_/B _07636_/B VGND VGND VPWR VPWR _07637_/B sky130_fd_sc_hd__or2_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07567_ _07578_/A _07578_/B VGND VGND VPWR VPWR _07567_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09306_ _13291_/Q _13529_/Q _09310_/S VGND VGND VPWR VPWR _09307_/A sky130_fd_sc_hd__mux2_1
X_06518_ _06499_/A _06499_/B _06499_/C _06517_/Y VGND VGND VPWR VPWR _06519_/B sky130_fd_sc_hd__o31ai_1
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07498_ _07498_/A _07498_/B _07504_/D VGND VGND VPWR VPWR _07498_/Y sky130_fd_sc_hd__nand3_1
XFILLER_10_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09237_ _13546_/Q _09237_/B VGND VGND VPWR VPWR _09241_/B sky130_fd_sc_hd__xor2_1
X_06449_ _06449_/A _06449_/B VGND VGND VPWR VPWR _06452_/A sky130_fd_sc_hd__or2_1
XFILLER_10_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09168_ _09106_/X _09173_/B _09167_/Y _07426_/X VGND VGND VPWR VPWR _13535_/D sky130_fd_sc_hd__a31o_1
XFILLER_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08119_ _08164_/A _13354_/Q _08119_/C VGND VGND VPWR VPWR _08123_/A sky130_fd_sc_hd__and3_1
X_09099_ _09099_/A _09099_/B _13526_/Q VGND VGND VPWR VPWR _09099_/X sky130_fd_sc_hd__or3b_1
X_11130_ _11130_/A VGND VGND VPWR VPWR _11130_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11061_ _11106_/A _11061_/B VGND VGND VPWR VPWR _11061_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10012_ _10095_/S VGND VGND VPWR VPWR _14048_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11963_ _14298_/Q _11962_/X _11966_/S VGND VGND VPWR VPWR _11964_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_83_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _14588_/CLK sky130_fd_sc_hd__clkbuf_16
X_13702_ _13702_/CLK _13702_/D VGND VGND VPWR VPWR hold508/A sky130_fd_sc_hd__dfxtp_1
X_10914_ _10914_/A VGND VGND VPWR VPWR _10914_/X sky130_fd_sc_hd__buf_2
X_14682_ _14688_/CLK hold278/X VGND VGND VPWR VPWR _14682_/Q sky130_fd_sc_hd__dfxtp_1
X_11894_ _14244_/Q _11522_/X _11894_/S VGND VGND VPWR VPWR _11895_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13633_ _13855_/CLK hold300/X VGND VGND VPWR VPWR _13633_/Q sky130_fd_sc_hd__dfxtp_1
X_10845_ _10845_/A VGND VGND VPWR VPWR _13182_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13564_ _13574_/CLK hold380/X VGND VGND VPWR VPWR _13564_/Q sky130_fd_sc_hd__dfxtp_1
X_10776_ _10776_/A VGND VGND VPWR VPWR _13051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12515_ _11285_/X _14704_/Q _12521_/S VGND VGND VPWR VPWR _12516_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13495_ _13704_/CLK hold110/X VGND VGND VPWR VPWR _13495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12446_ _14655_/Q _14701_/Q _12450_/S VGND VGND VPWR VPWR _12447_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12377_ _12377_/A VGND VGND VPWR VPWR _12386_/S sky130_fd_sc_hd__buf_2
XFILLER_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14116_ _14605_/CLK hold27/X VGND VGND VPWR VPWR hold428/A sky130_fd_sc_hd__dfxtp_1
X_11328_ _11328_/A VGND VGND VPWR VPWR _13769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14047_ _14047_/CLK hold355/X VGND VGND VPWR VPWR _14047_/Q sky130_fd_sc_hd__dfxtp_1
X_11259_ _14619_/Q _14581_/Q _14512_/Q _14464_/Q _12586_/A _11092_/A VGND VGND VPWR
+ VPWR _11260_/A sky130_fd_sc_hd__mux4_1
XFILLER_68_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_74_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _13593_/CLK sky130_fd_sc_hd__clkbuf_16
X_08470_ _08470_/A VGND VGND VPWR VPWR _08645_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07421_ _07400_/A _07418_/X _07435_/A VGND VGND VPWR VPWR _09164_/B sky130_fd_sc_hd__o21a_1
XFILLER_90_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07352_ _07364_/A _07359_/C VGND VGND VPWR VPWR _09126_/B sky130_fd_sc_hd__and2_2
XFILLER_149_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06303_ _13872_/Q _13856_/Q _06313_/S VGND VGND VPWR VPWR _06304_/A sky130_fd_sc_hd__mux2_1
X_07283_ _07231_/Y _07400_/B _07282_/X _07228_/X VGND VGND VPWR VPWR _07283_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09022_ _09022_/A VGND VGND VPWR VPWR _12747_/D sky130_fd_sc_hd__clkbuf_1
X_06234_ _06245_/B VGND VGND VPWR VPWR _12036_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold200 hold200/A VGND VGND VPWR VPWR hold200/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06165_ _13856_/Q _11836_/B VGND VGND VPWR VPWR _06166_/A sky130_fd_sc_hd__and2_1
Xhold211 hold211/A VGND VGND VPWR VPWR hold211/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold222 hold222/A VGND VGND VPWR VPWR hold222/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold233 hold233/A VGND VGND VPWR VPWR hold233/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold244 hold244/A VGND VGND VPWR VPWR hold244/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold255 hold255/A VGND VGND VPWR VPWR hold255/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06096_ _06096_/A VGND VGND VPWR VPWR _13938_/D sky130_fd_sc_hd__clkbuf_1
Xhold266 hold266/A VGND VGND VPWR VPWR hold266/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold277 hold277/A VGND VGND VPWR VPWR hold277/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold288 hold288/A VGND VGND VPWR VPWR hold288/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold299 hold299/A VGND VGND VPWR VPWR hold299/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09924_ _13487_/Q _13676_/Q _09924_/S VGND VGND VPWR VPWR _09925_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09855_ _09855_/A VGND VGND VPWR VPWR _09855_/X sky130_fd_sc_hd__buf_2
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08806_ _08828_/A _08819_/A _08833_/C VGND VGND VPWR VPWR _08826_/A sky130_fd_sc_hd__and3_1
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06998_ _13028_/Q _08015_/B VGND VGND VPWR VPWR _06999_/B sky130_fd_sc_hd__nor2_1
X_09786_ _09776_/X _09783_/Y _09785_/Y VGND VGND VPWR VPWR _13676_/D sky130_fd_sc_hd__a21oi_1
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05949_ _13867_/Q _13868_/Q _13869_/Q _13870_/Q VGND VGND VPWR VPWR _05950_/C sky130_fd_sc_hd__and4_1
X_08737_ _13458_/Q _08746_/A VGND VGND VPWR VPWR _08739_/C sky130_fd_sc_hd__xor2_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_65_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _13534_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _13449_/Q _09464_/B _08662_/A VGND VGND VPWR VPWR _08668_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07619_ _07791_/A VGND VGND VPWR VPWR _07738_/A sky130_fd_sc_hd__buf_2
XFILLER_41_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ _13443_/Q _08577_/B _08587_/A VGND VGND VPWR VPWR _08621_/B sky130_fd_sc_hd__a21oi_1
XFILLER_42_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10630_ _14523_/Q _14522_/Q _14525_/Q _14524_/Q VGND VGND VPWR VPWR _10630_/X sky130_fd_sc_hd__or4_1
X_10561_ _10562_/A _10562_/B _10562_/C VGND VGND VPWR VPWR _10570_/B sky130_fd_sc_hd__o21ai_1
XFILLER_128_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12300_ _14566_/Q _11978_/X _12302_/S VGND VGND VPWR VPWR _12301_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13280_ _13280_/CLK _13280_/D repeater59/X VGND VGND VPWR VPWR _13280_/Q sky130_fd_sc_hd__dfrtp_1
X_10492_ _10492_/A VGND VGND VPWR VPWR _14010_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12231_ _11285_/X _14532_/Q _12237_/S VGND VGND VPWR VPWR _12232_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12162_ _12162_/A VGND VGND VPWR VPWR _14493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11113_ _11065_/X _11110_/X _11112_/X _11086_/X VGND VGND VPWR VPWR _11113_/X sky130_fd_sc_hd__o211a_1
X_12093_ _11375_/X _14464_/Q _12093_/S VGND VGND VPWR VPWR _12094_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11044_ _11186_/A VGND VGND VPWR VPWR _11044_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_56_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _14645_/CLK sky130_fd_sc_hd__clkbuf_16
X_12995_ _14636_/CLK hold211/X VGND VGND VPWR VPWR hold159/A sky130_fd_sc_hd__dfxtp_4
XFILLER_17_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14734_ _14749_/CLK _14734_/D VGND VGND VPWR VPWR _14734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11946_ _14279_/Q _11519_/X _11948_/S VGND VGND VPWR VPWR _11947_/A sky130_fd_sc_hd__mux2_1
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14665_ _14720_/CLK _14665_/D VGND VGND VPWR VPWR _14665_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _11877_/A VGND VGND VPWR VPWR _11886_/S sky130_fd_sc_hd__buf_2
XFILLER_32_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13616_ _13617_/CLK _13616_/D repeater57/X VGND VGND VPWR VPWR _13616_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10828_ _10828_/A VGND VGND VPWR VPWR _13175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14596_ _14749_/CLK _14596_/D VGND VGND VPWR VPWR _14596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13547_ _14082_/CLK _13547_/D _12609_/A VGND VGND VPWR VPWR _13547_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_158_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10759_ _10781_/A VGND VGND VPWR VPWR _10768_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13478_ _14250_/CLK hold209/X VGND VGND VPWR VPWR _13478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12429_ _12463_/A VGND VGND VPWR VPWR _12480_/S sky130_fd_sc_hd__buf_2
XFILLER_126_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07970_ _07970_/A _07970_/B _07970_/C VGND VGND VPWR VPWR _07970_/X sky130_fd_sc_hd__or3_1
XFILLER_87_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06921_ _13018_/Q _06938_/B VGND VGND VPWR VPWR _06932_/A sky130_fd_sc_hd__and2_1
XFILLER_110_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09640_ _13416_/Q _13614_/Q _09642_/S VGND VGND VPWR VPWR _09641_/A sky130_fd_sc_hd__mux2_1
X_06852_ _06852_/A _06852_/B VGND VGND VPWR VPWR _06852_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09571_ _09568_/Y _09569_/X _09564_/A _09565_/Y VGND VGND VPWR VPWR _09571_/X sky130_fd_sc_hd__a211o_1
X_06783_ _06841_/B _06645_/X _06783_/S VGND VGND VPWR VPWR _06783_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_47_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _14432_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08522_ _08532_/B _08536_/A VGND VGND VPWR VPWR _08523_/A sky130_fd_sc_hd__and2_1
XFILLER_36_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08453_ _08671_/B _08450_/C _08450_/D _08671_/A VGND VGND VPWR VPWR _09367_/C sky130_fd_sc_hd__a22o_1
XFILLER_51_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07404_ _13142_/Q _09153_/B _09153_/C VGND VGND VPWR VPWR _07414_/B sky130_fd_sc_hd__and3_1
X_08384_ _13089_/Q _13370_/Q _08384_/S VGND VGND VPWR VPWR _08385_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07335_ _07335_/A _07349_/B VGND VGND VPWR VPWR _09118_/B sky130_fd_sc_hd__xnor2_2
XFILLER_149_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07266_ _07266_/A VGND VGND VPWR VPWR _07428_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09005_ _09005_/A VGND VGND VPWR VPWR _14255_/D sky130_fd_sc_hd__clkbuf_1
X_06217_ _06324_/A _06324_/B _06216_/Y VGND VGND VPWR VPWR _06322_/S sky130_fd_sc_hd__a21oi_1
XFILLER_136_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07197_ _07197_/A _07197_/B VGND VGND VPWR VPWR _07198_/B sky130_fd_sc_hd__or2_1
XFILLER_105_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06148_ _06290_/S VGND VGND VPWR VPWR _10121_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_144_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06079_ _10034_/S VGND VGND VPWR VPWR _13965_/D sky130_fd_sc_hd__inv_2
XFILLER_59_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09907_ _13479_/Q _13668_/Q _09913_/S VGND VGND VPWR VPWR _09908_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09838_ _13682_/Q _09838_/B VGND VGND VPWR VPWR _09839_/B sky130_fd_sc_hd__nor2_1
XFILLER_47_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09769_ _13675_/Q _09769_/B VGND VGND VPWR VPWR _09770_/B sky130_fd_sc_hd__nor2_1
XFILLER_73_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _13263_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11800_ _13571_/Q _11806_/B VGND VGND VPWR VPWR _11801_/A sky130_fd_sc_hd__and2_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12780_ _13565_/CLK _12780_/D VGND VGND VPWR VPWR hold374/A sky130_fd_sc_hd__dfxtp_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _11731_/A VGND VGND VPWR VPWR _14057_/D sky130_fd_sc_hd__clkbuf_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14450_ _14712_/CLK _14450_/D VGND VGND VPWR VPWR _14450_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _11662_/A VGND VGND VPWR VPWR _14014_/D sky130_fd_sc_hd__clkbuf_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13401_ _13596_/CLK hold460/X VGND VGND VPWR VPWR _13401_/Q sky130_fd_sc_hd__dfxtp_1
X_10613_ _14281_/Q _14291_/Q VGND VGND VPWR VPWR _10613_/X sky130_fd_sc_hd__and2_1
XFILLER_41_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14381_ _14397_/CLK hold296/X VGND VGND VPWR VPWR hold230/A sky130_fd_sc_hd__dfxtp_1
X_11593_ _12680_/Q _11593_/B VGND VGND VPWR VPWR _11594_/A sky130_fd_sc_hd__and2_1
XFILLER_6_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10544_ _10567_/A _12990_/D _10557_/B _10509_/A VGND VGND VPWR VPWR _10545_/A sky130_fd_sc_hd__a22o_1
X_13332_ _14605_/CLK _13332_/D VGND VGND VPWR VPWR _13332_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10475_ _10485_/A _10485_/B _10456_/C _10474_/Y VGND VGND VPWR VPWR _10476_/B sky130_fd_sc_hd__a31o_1
X_13263_ _13263_/CLK _13263_/D hold1/X VGND VGND VPWR VPWR _13263_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12214_ _12214_/A _12214_/B VGND VGND VPWR VPWR _14515_/D sky130_fd_sc_hd__nor2_1
X_13194_ _13606_/CLK _13194_/D VGND VGND VPWR VPWR hold521/A sky130_fd_sc_hd__dfxtp_1
XFILLER_163_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12145_ _14487_/Q _12022_/X _12147_/S VGND VGND VPWR VPWR _12146_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12076_ _12076_/A VGND VGND VPWR VPWR _12085_/S sky130_fd_sc_hd__buf_2
XFILLER_77_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11027_ _13323_/Q _11008_/X _11016_/X _11026_/Y VGND VGND VPWR VPWR _13323_/D sky130_fd_sc_hd__o22a_1
XFILLER_77_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _13298_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12978_ _13280_/CLK hold256/X VGND VGND VPWR VPWR _12978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14717_ _14717_/CLK _14717_/D VGND VGND VPWR VPWR _14717_/Q sky130_fd_sc_hd__dfxtp_1
X_11929_ _14271_/Q _11494_/X _11929_/S VGND VGND VPWR VPWR _11930_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14648_ _14703_/CLK _14648_/D VGND VGND VPWR VPWR _14648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_17 input26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 _13318_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14579_ _14579_/CLK _14579_/D VGND VGND VPWR VPWR _14579_/Q sky130_fd_sc_hd__dfxtp_1
X_07120_ _07120_/A _07150_/A VGND VGND VPWR VPWR _07121_/B sky130_fd_sc_hd__nor2_1
XFILLER_146_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07051_ _07058_/B _07051_/B VGND VGND VPWR VPWR _07053_/B sky130_fd_sc_hd__xnor2_1
XFILLER_146_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06002_ hold173/A _13564_/Q _06002_/C _06002_/D VGND VGND VPWR VPWR _06002_/Y sky130_fd_sc_hd__nor4_2
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07953_ _07972_/A _07953_/B VGND VGND VPWR VPWR _07953_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06904_ _06914_/A _06904_/B VGND VGND VPWR VPWR _06924_/B sky130_fd_sc_hd__nand2_1
X_07884_ _07885_/D _07892_/B _07884_/C _07892_/D VGND VGND VPWR VPWR _07884_/X sky130_fd_sc_hd__or4_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09623_ _13408_/Q _13606_/Q _09631_/S VGND VGND VPWR VPWR _09624_/A sky130_fd_sc_hd__mux2_1
X_06835_ _06824_/X _06826_/X _06828_/X _06834_/Y VGND VGND VPWR VPWR _06846_/B sky130_fd_sc_hd__a31o_1
XFILLER_55_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09554_ _09502_/X _09556_/B _09553_/Y _09506_/X VGND VGND VPWR VPWR _13615_/D sky130_fd_sc_hd__a31o_1
XFILLER_83_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06766_ _06766_/A VGND VGND VPWR VPWR _13005_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08505_ _14255_/Q _14253_/Q _08506_/S VGND VGND VPWR VPWR _08505_/X sky130_fd_sc_hd__mux2_1
X_09485_ _09510_/A _09509_/A VGND VGND VPWR VPWR _09485_/X sky130_fd_sc_hd__or2_1
X_06697_ _06712_/A _06696_/Y VGND VGND VPWR VPWR _06700_/A sky130_fd_sc_hd__or2b_1
XFILLER_62_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08436_ _08671_/B _08450_/C VGND VGND VPWR VPWR _09370_/B sky130_fd_sc_hd__xor2_4
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08367_ _13081_/Q _13362_/Q _08373_/S VGND VGND VPWR VPWR _08368_/A sky130_fd_sc_hd__mux2_1
X_07318_ _07318_/A _07318_/B VGND VGND VPWR VPWR _07322_/A sky130_fd_sc_hd__or2_1
X_08298_ _09116_/S VGND VGND VPWR VPWR _08298_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07249_ _07311_/A _07461_/B _07249_/C _07249_/D VGND VGND VPWR VPWR _09086_/B sky130_fd_sc_hd__nand4_4
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10260_ _10251_/X _10259_/X _14556_/D VGND VGND VPWR VPWR _10260_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10191_ _10226_/A _14362_/Q VGND VGND VPWR VPWR _10230_/A sky130_fd_sc_hd__xnor2_1
XFILLER_105_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13950_ _13964_/CLK _13950_/D VGND VGND VPWR VPWR _13950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12901_ _13274_/CLK _12901_/D hold1/X VGND VGND VPWR VPWR _12901_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13881_ _14657_/CLK hold236/X VGND VGND VPWR VPWR hold427/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _14327_/CLK _12832_/D VGND VGND VPWR VPWR hold430/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _13700_/CLK _12763_/D VGND VGND VPWR VPWR hold202/A sky130_fd_sc_hd__dfxtp_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _14610_/CLK _14502_/D VGND VGND VPWR VPWR _14502_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _12619_/A _12041_/C _12621_/A VGND VGND VPWR VPWR _11749_/A sky130_fd_sc_hd__nand3b_4
XFILLER_42_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _13304_/CLK _12694_/D VGND VGND VPWR VPWR hold105/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _14435_/CLK _14433_/D VGND VGND VPWR VPWR _14433_/Q sky130_fd_sc_hd__dfxtp_1
X_11645_ _13998_/Q _11510_/X _11645_/S VGND VGND VPWR VPWR _11646_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput15 data_i[22] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__buf_6
X_14364_ _14557_/CLK hold497/X VGND VGND VPWR VPWR hold304/A sky130_fd_sc_hd__dfxtp_1
Xinput26 data_i[9] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_4
X_11576_ _11576_/A VGND VGND VPWR VPWR _11585_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_155_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13315_ _14108_/CLK hold290/X VGND VGND VPWR VPWR _13315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10527_ _13815_/Q VGND VGND VPWR VPWR _10557_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14295_ _14742_/CLK _14295_/D VGND VGND VPWR VPWR _14295_/Q sky130_fd_sc_hd__dfxtp_1
X_13246_ _14687_/CLK _13246_/D VGND VGND VPWR VPWR _13518_/D sky130_fd_sc_hd__dfxtp_2
X_10458_ hold79/A _10465_/A VGND VGND VPWR VPWR _10476_/A sky130_fd_sc_hd__and2_1
XFILLER_143_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10389_ _10390_/A _10390_/B VGND VGND VPWR VPWR _10407_/A sky130_fd_sc_hd__and2_1
XFILLER_97_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13177_ _13596_/CLK _13177_/D VGND VGND VPWR VPWR hold75/A sky130_fd_sc_hd__dfxtp_1
XFILLER_151_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12128_ _14479_/Q _11997_/X _12128_/S VGND VGND VPWR VPWR _12129_/A sky130_fd_sc_hd__mux2_1
X_12059_ _11304_/X _14448_/Q _12063_/S VGND VGND VPWR VPWR _12060_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06620_ _12903_/Q _06620_/B _06620_/C VGND VGND VPWR VPWR _06620_/X sky130_fd_sc_hd__and3_1
XFILLER_65_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06551_ _12910_/Q VGND VGND VPWR VPWR _06609_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_33_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09270_ _13551_/Q _09270_/B VGND VGND VPWR VPWR _09272_/A sky130_fd_sc_hd__and2_1
X_06482_ _06482_/A VGND VGND VPWR VPWR _06502_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08221_ _13363_/Q _08226_/B VGND VGND VPWR VPWR _08234_/A sky130_fd_sc_hd__nor2_1
X_08152_ _08220_/B _13356_/Q _08152_/C VGND VGND VPWR VPWR _08152_/X sky130_fd_sc_hd__and3_1
X_07103_ _07218_/S VGND VGND VPWR VPWR _07199_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_119_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08083_ _08083_/A VGND VGND VPWR VPWR _12701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_9_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _13274_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_162_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07034_ _13036_/D _07034_/B VGND VGND VPWR VPWR _07034_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_134_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08985_ _08985_/A _08985_/B VGND VGND VPWR VPWR _08986_/B sky130_fd_sc_hd__or2_1
XFILLER_87_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07936_ _13270_/Q _07947_/B VGND VGND VPWR VPWR _07937_/B sky130_fd_sc_hd__or2_1
XFILLER_130_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07867_ _07885_/C _07892_/A _07866_/X VGND VGND VPWR VPWR _07867_/Y sky130_fd_sc_hd__o21ai_1
X_09606_ _09606_/A VGND VGND VPWR VPWR _12817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06818_ _06825_/B _06825_/C VGND VGND VPWR VPWR _06820_/C sky130_fd_sc_hd__or2_1
X_07798_ _07791_/Y _07797_/Y _07800_/S VGND VGND VPWR VPWR _07799_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09537_ _09510_/A _09535_/X _09536_/Y _09508_/Y VGND VGND VPWR VPWR _09548_/A sky130_fd_sc_hd__o211ai_4
XFILLER_25_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06749_ _13039_/Q VGND VGND VPWR VPWR _06782_/A sky130_fd_sc_hd__inv_2
X_09468_ _09477_/A _09468_/B VGND VGND VPWR VPWR _09475_/B sky130_fd_sc_hd__or2_1
XFILLER_24_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08419_ _08419_/A VGND VGND VPWR VPWR _12740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09399_ _13595_/Q _09399_/B VGND VGND VPWR VPWR _09419_/C sky130_fd_sc_hd__xnor2_4
X_11430_ _13737_/Q _11438_/B VGND VGND VPWR VPWR _11431_/A sky130_fd_sc_hd__and2_1
XFILLER_11_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11361_ _11361_/A VGND VGND VPWR VPWR _13775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13100_ _14555_/CLK hold392/X VGND VGND VPWR VPWR _13100_/Q sky130_fd_sc_hd__dfxtp_1
X_10312_ _10312_/A _10312_/B VGND VGND VPWR VPWR _13475_/D sky130_fd_sc_hd__xnor2_1
XFILLER_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11292_ _13758_/Q _11291_/X _11295_/S VGND VGND VPWR VPWR _11293_/A sky130_fd_sc_hd__mux2_1
X_14080_ _14082_/CLK _14080_/D VGND VGND VPWR VPWR _14080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10243_ _14523_/D _10242_/X _14557_/D VGND VGND VPWR VPWR _10244_/A sky130_fd_sc_hd__mux2_1
X_13031_ _13031_/CLK _13031_/D VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__dfxtp_1
XFILLER_106_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10174_ _10169_/X _10173_/X _14292_/D VGND VGND VPWR VPWR _10175_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13933_ _14179_/CLK hold370/X VGND VGND VPWR VPWR _13933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13864_ _14075_/CLK _13864_/D VGND VGND VPWR VPWR _13864_/Q sky130_fd_sc_hd__dfxtp_1
X_12815_ _13653_/CLK _12815_/D VGND VGND VPWR VPWR hold153/A sky130_fd_sc_hd__dfxtp_1
X_13795_ _13843_/CLK _13795_/D VGND VGND VPWR VPWR _13795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12746_ _13702_/CLK _12746_/D VGND VGND VPWR VPWR hold265/A sky130_fd_sc_hd__dfxtp_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12677_ _13296_/CLK _12677_/D VGND VGND VPWR VPWR hold338/A sky130_fd_sc_hd__dfxtp_1
XFILLER_147_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14416_ _14424_/CLK _14416_/D VGND VGND VPWR VPWR _14416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11628_ _13990_/Q _11485_/X _11634_/S VGND VGND VPWR VPWR _11629_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14347_ _14357_/CLK hold373/X VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__dfxtp_1
X_11559_ _13638_/Q _11563_/B VGND VGND VPWR VPWR _11560_/A sky130_fd_sc_hd__and2_1
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14278_ _14724_/CLK _14278_/D VGND VGND VPWR VPWR _14278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13229_ _13610_/CLK hold457/X VGND VGND VPWR VPWR _13229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05982_ _14095_/Q _14096_/Q _14097_/Q _14098_/Q VGND VGND VPWR VPWR _05983_/C sky130_fd_sc_hd__or4_1
X_08770_ _08770_/A _08770_/B VGND VGND VPWR VPWR _08770_/Y sky130_fd_sc_hd__nor2_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07721_ _07721_/A _07772_/D VGND VGND VPWR VPWR _07729_/A sky130_fd_sc_hd__nand2_1
XFILLER_111_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07652_ _07664_/A _07664_/B VGND VGND VPWR VPWR _07654_/B sky130_fd_sc_hd__xnor2_1
XFILLER_19_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06603_ _12900_/Q _06607_/D _06599_/X VGND VGND VPWR VPWR _06604_/B sky130_fd_sc_hd__o21ai_1
XFILLER_53_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07583_ _07583_/A _07583_/B _07583_/C VGND VGND VPWR VPWR _07583_/Y sky130_fd_sc_hd__nand3_1
XFILLER_40_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09322_ _09322_/A VGND VGND VPWR VPWR _12788_/D sky130_fd_sc_hd__clkbuf_1
X_06534_ _12888_/Q _06534_/B VGND VGND VPWR VPWR _06535_/B sky130_fd_sc_hd__nor2_1
XFILLER_22_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09253_ _09125_/X _09252_/X _07486_/X VGND VGND VPWR VPWR _13548_/D sky130_fd_sc_hd__a21o_1
X_06465_ _06465_/A _06465_/B VGND VGND VPWR VPWR _06465_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_21_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08204_ _08204_/A _08204_/B VGND VGND VPWR VPWR _08204_/Y sky130_fd_sc_hd__xnor2_1
X_09184_ _13538_/Q _09188_/B VGND VGND VPWR VPWR _09189_/B sky130_fd_sc_hd__xnor2_1
XFILLER_21_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06396_ _10346_/A _06504_/B _06395_/X _06429_/B VGND VGND VPWR VPWR _06405_/B sky130_fd_sc_hd__a22o_1
X_08135_ _13356_/Q _08135_/B VGND VGND VPWR VPWR _08136_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08066_ _08066_/A VGND VGND VPWR VPWR _12693_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07017_ hold425/A _07063_/B VGND VGND VPWR VPWR _07045_/C sky130_fd_sc_hd__and2_1
XFILLER_1_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08968_ _08984_/A _08968_/B VGND VGND VPWR VPWR _08970_/C sky130_fd_sc_hd__nand2_1
XFILLER_29_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07919_ _13267_/Q _07911_/B _07917_/B _07918_/Y VGND VGND VPWR VPWR _07919_/Y sky130_fd_sc_hd__a22oi_1
X_08899_ _08899_/A _08899_/B VGND VGND VPWR VPWR _08901_/A sky130_fd_sc_hd__nor2_1
XFILLER_56_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10930_ _12645_/A _10919_/X _10926_/X _10929_/X VGND VGND VPWR VPWR _10930_/X sky130_fd_sc_hd__o211a_1
XFILLER_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10861_ _13148_/Q _10863_/B VGND VGND VPWR VPWR _10862_/A sky130_fd_sc_hd__and2_1
X_12600_ _12604_/C _12599_/Y _12580_/X VGND VGND VPWR VPWR _14730_/D sky130_fd_sc_hd__o21ai_1
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13580_ _14275_/CLK hold349/X VGND VGND VPWR VPWR _13580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10792_ _10803_/A VGND VGND VPWR VPWR _10801_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12531_ _12531_/A VGND VGND VPWR VPWR _14711_/D sky130_fd_sc_hd__clkbuf_1
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12462_ _12462_/A VGND VGND VPWR VPWR _14662_/D sky130_fd_sc_hd__clkbuf_1
X_14201_ _14201_/CLK _14201_/D VGND VGND VPWR VPWR _14201_/Q sky130_fd_sc_hd__dfxtp_1
X_11413_ _11413_/A VGND VGND VPWR VPWR _13798_/D sky130_fd_sc_hd__clkbuf_1
X_12393_ _12393_/A VGND VGND VPWR VPWR _14618_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14132_ _14716_/CLK hold330/X VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__dfxtp_1
X_11344_ _13772_/Q _11343_/X _11355_/S VGND VGND VPWR VPWR _11345_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14063_ _14543_/CLK _14063_/D VGND VGND VPWR VPWR _14063_/Q sky130_fd_sc_hd__dfxtp_1
X_11275_ _12662_/D _12661_/D _12662_/Q _11274_/Y VGND VGND VPWR VPWR _12582_/A sky130_fd_sc_hd__o31ai_4
XFILLER_79_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13014_ _13304_/CLK _13014_/D repeater59/X VGND VGND VPWR VPWR _13014_/Q sky130_fd_sc_hd__dfrtp_1
X_10226_ _10226_/A _14377_/Q VGND VGND VPWR VPWR _10236_/B sky130_fd_sc_hd__xnor2_1
XFILLER_79_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10157_ _10157_/A VGND VGND VPWR VPWR _14288_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_10088_ _10088_/A VGND VGND VPWR VPWR _13904_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13916_ _13978_/CLK _13916_/D VGND VGND VPWR VPWR hold160/A sky130_fd_sc_hd__dfxtp_1
XFILLER_90_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13847_ _14180_/CLK _13847_/D VGND VGND VPWR VPWR _13847_/Q sky130_fd_sc_hd__dfxtp_1
X_13778_ _14726_/CLK _13778_/D VGND VGND VPWR VPWR _13778_/Q sky130_fd_sc_hd__dfxtp_1
X_12729_ _13617_/CLK _12729_/D VGND VGND VPWR VPWR hold424/A sky130_fd_sc_hd__dfxtp_1
X_06250_ _14079_/Q _14080_/Q _14081_/Q _14082_/Q VGND VGND VPWR VPWR _06250_/X sky130_fd_sc_hd__or4_1
XFILLER_164_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06181_ _06179_/X _06180_/X _11836_/B VGND VGND VPWR VPWR _14196_/D sky130_fd_sc_hd__o21a_1
XFILLER_144_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold404 hold404/A VGND VGND VPWR VPWR hold404/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold415 hold415/A VGND VGND VPWR VPWR hold415/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold426 hold426/A VGND VGND VPWR VPWR hold426/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold437 hold437/A VGND VGND VPWR VPWR hold437/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold448 hold448/A VGND VGND VPWR VPWR hold448/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09940_ _13494_/Q _13683_/Q _09946_/S VGND VGND VPWR VPWR _09941_/A sky130_fd_sc_hd__mux2_1
Xhold459 hold459/A VGND VGND VPWR VPWR hold459/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_143_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _13689_/Q _09868_/A _09776_/X VGND VGND VPWR VPWR _09872_/B sky130_fd_sc_hd__o21ai_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08822_ _13473_/D _08822_/B VGND VGND VPWR VPWR _08822_/Y sky130_fd_sc_hd__xnor2_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08753_ _13459_/Q _09581_/B _08758_/A _08757_/A VGND VGND VPWR VPWR _08754_/B sky130_fd_sc_hd__a22o_1
X_05965_ _13625_/Q _13626_/Q _13627_/Q _13628_/Q VGND VGND VPWR VPWR _05965_/X sky130_fd_sc_hd__and4_1
X_07704_ _07705_/A _07705_/B _07705_/C VGND VGND VPWR VPWR _07733_/A sky130_fd_sc_hd__a21o_1
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ _09493_/A VGND VGND VPWR VPWR _08684_/X sky130_fd_sc_hd__clkbuf_2
X_05896_ _13780_/Q VGND VGND VPWR VPWR hold516/A sky130_fd_sc_hd__clkinv_2
XFILLER_53_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07635_ _07635_/A _07635_/B VGND VGND VPWR VPWR _07636_/B sky130_fd_sc_hd__nor2_1
XFILLER_26_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07566_ _07566_/A _07566_/B VGND VGND VPWR VPWR _07578_/B sky130_fd_sc_hd__or2_1
XFILLER_53_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09305_ _09305_/A VGND VGND VPWR VPWR _12780_/D sky130_fd_sc_hd__clkbuf_1
X_06517_ _12884_/Q _06500_/B _06506_/A VGND VGND VPWR VPWR _06517_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07497_ _07498_/A _07498_/B _07504_/D VGND VGND VPWR VPWR _07497_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09236_ _09182_/X _09234_/Y _09235_/X _09215_/X VGND VGND VPWR VPWR _13545_/D sky130_fd_sc_hd__a31o_1
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06448_ _12880_/Q _06448_/B VGND VGND VPWR VPWR _06449_/B sky130_fd_sc_hd__nor2_1
XFILLER_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09167_ _09149_/B _09160_/B _09158_/X _09165_/Y VGND VGND VPWR VPWR _09167_/Y sky130_fd_sc_hd__o211ai_1
X_06379_ _13108_/D VGND VGND VPWR VPWR _06392_/A sky130_fd_sc_hd__inv_2
XFILLER_135_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08118_ _08114_/X _08116_/X _08220_/C _08208_/A VGND VGND VPWR VPWR _08120_/C sky130_fd_sc_hd__a2bb2o_1
XFILLER_163_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09098_ _13526_/Q _09098_/B VGND VGND VPWR VPWR _09109_/A sky130_fd_sc_hd__nor2_1
XFILLER_119_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08049_ _12962_/Q _13262_/Q _08051_/S VGND VGND VPWR VPWR _08050_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11060_ _14265_/Q _14656_/Q _13763_/Q _14711_/Q _11020_/X _11021_/X VGND VGND VPWR
+ VPWR _11061_/B sky130_fd_sc_hd__mux4_1
XFILLER_1_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10011_ _10052_/A _13910_/Q VGND VGND VPWR VPWR _10095_/S sky130_fd_sc_hd__xor2_2
XFILLER_77_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11962_ _14697_/Q VGND VGND VPWR VPWR _11962_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13701_ _13702_/CLK _13701_/D VGND VGND VPWR VPWR _13701_/Q sky130_fd_sc_hd__dfxtp_1
X_10913_ _12586_/A VGND VGND VPWR VPWR _10914_/A sky130_fd_sc_hd__buf_2
X_14681_ _14688_/CLK hold270/X VGND VGND VPWR VPWR _14681_/Q sky130_fd_sc_hd__dfxtp_1
X_11893_ _11893_/A VGND VGND VPWR VPWR _14243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13632_ _13855_/CLK hold409/X VGND VGND VPWR VPWR _13632_/Q sky130_fd_sc_hd__dfxtp_1
X_10844_ _13140_/Q _10852_/B VGND VGND VPWR VPWR _10845_/A sky130_fd_sc_hd__and2_1
XFILLER_71_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13563_ _13587_/CLK hold144/X VGND VGND VPWR VPWR _13563_/Q sky130_fd_sc_hd__dfxtp_1
X_10775_ _13009_/Q _10779_/B VGND VGND VPWR VPWR _10776_/A sky130_fd_sc_hd__and2_1
X_12514_ _12514_/A VGND VGND VPWR VPWR _14703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13494_ _13602_/CLK hold242/X VGND VGND VPWR VPWR _13494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12445_ _12445_/A VGND VGND VPWR VPWR _14654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12376_ _12376_/A VGND VGND VPWR VPWR _14610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14115_ _14605_/CLK hold428/X VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__dfxtp_1
XFILLER_141_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11327_ _13769_/Q _11326_/X _11327_/S VGND VGND VPWR VPWR _11328_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14046_ _14210_/CLK _14046_/D VGND VGND VPWR VPWR hold355/A sky130_fd_sc_hd__dfxtp_1
X_11258_ _11207_/X _11255_/X _11257_/X _12647_/A VGND VGND VPWR VPWR _11258_/X sky130_fd_sc_hd__o211a_1
XFILLER_141_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10209_ _10209_/A VGND VGND VPWR VPWR _14420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11189_ _11189_/A VGND VGND VPWR VPWR _11189_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07420_ _07420_/A VGND VGND VPWR VPWR _07435_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07351_ _07350_/A _07349_/A _07349_/B _07349_/C VGND VGND VPWR VPWR _07359_/C sky130_fd_sc_hd__a31o_1
XFILLER_148_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06302_ _06302_/A VGND VGND VPWR VPWR _14185_/D sky130_fd_sc_hd__clkbuf_1
X_07282_ _13660_/Q _13656_/Q _13658_/Q _13390_/Q _07247_/X _07267_/S VGND VGND VPWR
+ VPWR _07282_/X sky130_fd_sc_hd__mux4_1
X_06233_ _06233_/A VGND VGND VPWR VPWR _14386_/D sky130_fd_sc_hd__clkbuf_1
X_09021_ _13211_/Q _13440_/Q _09029_/S VGND VGND VPWR VPWR _09022_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06164_ _06175_/B VGND VGND VPWR VPWR _11836_/B sky130_fd_sc_hd__clkbuf_1
Xhold201 hold201/A VGND VGND VPWR VPWR hold201/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold212 hold212/A VGND VGND VPWR VPWR hold212/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold223 hold223/A VGND VGND VPWR VPWR hold223/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold234 hold234/A VGND VGND VPWR VPWR hold234/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_160_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06095_ _13792_/Q _11593_/B VGND VGND VPWR VPWR _06096_/A sky130_fd_sc_hd__and2_1
Xhold245 hold245/A VGND VGND VPWR VPWR hold245/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold256 hold256/A VGND VGND VPWR VPWR hold256/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold267 hold267/A VGND VGND VPWR VPWR hold267/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold278 hold278/A VGND VGND VPWR VPWR hold278/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09923_ _09923_/A VGND VGND VPWR VPWR _12849_/D sky130_fd_sc_hd__clkbuf_1
Xhold289 hold289/A VGND VGND VPWR VPWR hold289/X sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09854_ _09854_/A VGND VGND VPWR VPWR _13684_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08805_ _13516_/D _08851_/B VGND VGND VPWR VPWR _08833_/C sky130_fd_sc_hd__and2_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _09894_/A _09785_/B VGND VGND VPWR VPWR _09785_/Y sky130_fd_sc_hd__nor2_1
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06997_ _13028_/Q _08015_/B VGND VGND VPWR VPWR _06999_/A sky130_fd_sc_hd__and2_1
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08736_ _08739_/B _08734_/X _08735_/X VGND VGND VPWR VPWR _13457_/D sky130_fd_sc_hd__o21bai_1
X_05948_ _13871_/Q _13872_/Q _13873_/Q _13874_/Q VGND VGND VPWR VPWR _05950_/B sky130_fd_sc_hd__and4_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08667_ _13447_/Q _09450_/B _08644_/A VGND VGND VPWR VPWR _08667_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ _07618_/A VGND VGND VPWR VPWR _13656_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08598_ _13445_/Q _08602_/A VGND VGND VPWR VPWR _08620_/A sky130_fd_sc_hd__xnor2_1
XFILLER_41_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07549_ _13157_/Q _09270_/B VGND VGND VPWR VPWR _07556_/A sky130_fd_sc_hd__nand2_1
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10560_ _10565_/A _10560_/B VGND VGND VPWR VPWR _10562_/C sky130_fd_sc_hd__xnor2_1
X_09219_ _09226_/A _09219_/B VGND VGND VPWR VPWR _09242_/A sky130_fd_sc_hd__or2_1
X_10491_ _10498_/B _10491_/B VGND VGND VPWR VPWR _10492_/A sky130_fd_sc_hd__and2_1
X_12230_ _12230_/A VGND VGND VPWR VPWR _14531_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12161_ _14493_/Q _11965_/X _12161_/S VGND VGND VPWR VPWR _12162_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11112_ _11112_/A _11084_/X VGND VGND VPWR VPWR _11112_/X sky130_fd_sc_hd__or2b_1
XFILLER_1_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12092_ _12092_/A VGND VGND VPWR VPWR _14463_/D sky130_fd_sc_hd__clkbuf_1
X_11043_ _12649_/B VGND VGND VPWR VPWR _11108_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_3_0_clk clkbuf_4_3_0_clk/A VGND VGND VPWR VPWR clkbuf_4_3_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12994_ _14645_/CLK hold123/X VGND VGND VPWR VPWR _13116_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_45_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14733_ _14733_/CLK _14733_/D VGND VGND VPWR VPWR _14733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11945_ _11945_/A VGND VGND VPWR VPWR _14278_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _14733_/CLK _14664_/D VGND VGND VPWR VPWR _14664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ _11876_/A VGND VGND VPWR VPWR _14235_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13615_ _13619_/CLK _13615_/D repeater57/X VGND VGND VPWR VPWR _13615_/Q sky130_fd_sc_hd__dfrtp_1
X_10827_ _13133_/Q _10893_/A VGND VGND VPWR VPWR _10828_/A sky130_fd_sc_hd__and2_1
X_14595_ _14702_/CLK _14595_/D VGND VGND VPWR VPWR _14595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13546_ _13587_/CLK _13546_/D _12609_/A VGND VGND VPWR VPWR _13546_/Q sky130_fd_sc_hd__dfrtp_2
X_10758_ _10758_/A VGND VGND VPWR VPWR _13043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13477_ _14012_/CLK _13477_/D VGND VGND VPWR VPWR _13477_/Q sky130_fd_sc_hd__dfxtp_1
X_10689_ _10748_/B VGND VGND VPWR VPWR _10698_/B sky130_fd_sc_hd__clkbuf_1
X_12428_ _12510_/A _12428_/B VGND VGND VPWR VPWR _12463_/A sky130_fd_sc_hd__nor2_8
XFILLER_127_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12359_ _12359_/A VGND VGND VPWR VPWR _14602_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14029_ _14410_/CLK _14029_/D VGND VGND VPWR VPWR _14029_/Q sky130_fd_sc_hd__dfxtp_1
X_06920_ _06861_/X _06918_/X _06919_/Y _06907_/X VGND VGND VPWR VPWR _13017_/D sky130_fd_sc_hd__a31o_1
XFILLER_122_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06851_ _06851_/A _06851_/B VGND VGND VPWR VPWR _06858_/A sky130_fd_sc_hd__nor2_1
XFILLER_110_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09570_ _09564_/A _09565_/Y _09568_/Y _09569_/X VGND VGND VPWR VPWR _09570_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_67_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06782_ _06782_/A VGND VGND VPWR VPWR _06863_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08521_ _08521_/A _08552_/A VGND VGND VPWR VPWR _08536_/A sky130_fd_sc_hd__nand2_2
XFILLER_36_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08452_ _08535_/A VGND VGND VPWR VPWR _08671_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07403_ _09139_/B _07401_/B _07401_/C _07389_/A VGND VGND VPWR VPWR _09153_/C sky130_fd_sc_hd__o22ai_4
XFILLER_149_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08383_ _08383_/A VGND VGND VPWR VPWR _12724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07334_ _07327_/X _07330_/X _07333_/X _07311_/A VGND VGND VPWR VPWR _07349_/B sky130_fd_sc_hd__o211a_1
XFILLER_164_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07265_ _07224_/A _13663_/Q _13665_/Q _13661_/Q _07247_/X _07267_/S VGND VGND VPWR
+ VPWR _07388_/B sky130_fd_sc_hd__mux4_2
XFILLER_118_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09004_ _08997_/Y _09003_/Y _09006_/S VGND VGND VPWR VPWR _09005_/A sky130_fd_sc_hd__mux2_1
X_06216_ _06216_/A _06216_/B VGND VGND VPWR VPWR _06216_/Y sky130_fd_sc_hd__nor2_1
XFILLER_164_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07196_ _07196_/A _07196_/B _07196_/C VGND VGND VPWR VPWR _07197_/B sky130_fd_sc_hd__and3_1
X_06147_ _06292_/A _06292_/B _06146_/Y VGND VGND VPWR VPWR _06290_/S sky130_fd_sc_hd__a21oi_1
XFILLER_105_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06078_ _06257_/S VGND VGND VPWR VPWR _10034_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_132_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09906_ _09906_/A VGND VGND VPWR VPWR _12841_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09837_ _13682_/Q _09838_/B VGND VGND VPWR VPWR _09839_/A sky130_fd_sc_hd__and2_1
XFILLER_47_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09768_ _13675_/Q _09768_/B _09809_/C VGND VGND VPWR VPWR _09770_/A sky130_fd_sc_hd__and3_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _08633_/X _08718_/X _08684_/X VGND VGND VPWR VPWR _13455_/D sky130_fd_sc_hd__a21o_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _09699_/A VGND VGND VPWR VPWR _13669_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _11301_/X _14057_/Q _11736_/S VGND VGND VPWR VPWR _11731_/A sky130_fd_sc_hd__mux2_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _14014_/Q _11453_/X _11667_/S VGND VGND VPWR VPWR _11662_/A sky130_fd_sc_hd__mux2_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13400_ _13596_/CLK hold53/X VGND VGND VPWR VPWR _13400_/Q sky130_fd_sc_hd__dfxtp_1
X_10612_ _14050_/Q _10610_/X _10611_/X _14049_/Q _14038_/Q VGND VGND VPWR VPWR _14045_/D
+ sky130_fd_sc_hd__a221o_1
X_14380_ _14397_/CLK _14380_/D VGND VGND VPWR VPWR hold296/A sky130_fd_sc_hd__dfxtp_1
X_11592_ _11592_/A VGND VGND VPWR VPWR _13877_/D sky130_fd_sc_hd__clkbuf_1
X_13331_ _14717_/CLK _13331_/D VGND VGND VPWR VPWR _13331_/Q sky130_fd_sc_hd__dfxtp_1
X_10543_ _10555_/B _10557_/A _10531_/B VGND VGND VPWR VPWR _10549_/B sky130_fd_sc_hd__o21ai_1
XFILLER_10_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13262_ _13263_/CLK _13262_/D hold1/X VGND VGND VPWR VPWR _13262_/Q sky130_fd_sc_hd__dfrtp_1
X_10474_ _10474_/A VGND VGND VPWR VPWR _10474_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12213_ _14122_/Q _12215_/C _12205_/X VGND VGND VPWR VPWR _12214_/B sky130_fd_sc_hd__o21ai_1
XFILLER_6_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13193_ _13605_/CLK _13193_/D VGND VGND VPWR VPWR hold246/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12144_ _12144_/A VGND VGND VPWR VPWR _14486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12075_ _12075_/A VGND VGND VPWR VPWR _14455_/D sky130_fd_sc_hd__clkbuf_1
X_11026_ _11037_/A _11026_/B VGND VGND VPWR VPWR _11026_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12977_ _13280_/CLK hold258/X VGND VGND VPWR VPWR _12977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11928_ _11928_/A VGND VGND VPWR VPWR _14270_/D sky130_fd_sc_hd__clkbuf_1
X_14716_ _14716_/CLK _14716_/D VGND VGND VPWR VPWR _14716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14647_ _14647_/CLK _14647_/D VGND VGND VPWR VPWR _14647_/Q sky130_fd_sc_hd__dfxtp_1
X_11859_ _11859_/A VGND VGND VPWR VPWR _14227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_18 input26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_29 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14578_ _14579_/CLK _14578_/D VGND VGND VPWR VPWR _14578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13529_ _13534_/CLK _13529_/D hold1/X VGND VGND VPWR VPWR _13529_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07050_ _07028_/B _07032_/B _07028_/A VGND VGND VPWR VPWR _07051_/B sky130_fd_sc_hd__o21ba_1
X_06001_ _13577_/Q _13578_/Q _13579_/Q _06001_/D VGND VGND VPWR VPWR _06002_/D sky130_fd_sc_hd__or4_1
XFILLER_161_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07952_ _07972_/A _07953_/B VGND VGND VPWR VPWR _07952_/X sky130_fd_sc_hd__or2_1
XFILLER_68_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06903_ _13015_/Q _07963_/B VGND VGND VPWR VPWR _06904_/B sky130_fd_sc_hd__or2_1
XFILLER_68_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07883_ _07881_/A _07886_/C _07886_/D VGND VGND VPWR VPWR _07893_/B sky130_fd_sc_hd__o21ba_1
XFILLER_29_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09622_ _09644_/A VGND VGND VPWR VPWR _09631_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_68_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06834_ _06846_/A _06834_/B VGND VGND VPWR VPWR _06834_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09553_ _09559_/A _09553_/B _09553_/C VGND VGND VPWR VPWR _09553_/Y sky130_fd_sc_hd__nand3_1
X_06765_ _06757_/B _06762_/Y _07843_/S VGND VGND VPWR VPWR _06766_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08504_ _09365_/A VGND VGND VPWR VPWR _08504_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_70_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09484_ _09484_/A _09484_/B VGND VGND VPWR VPWR _09509_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06696_ _06719_/A _06696_/B _13001_/Q VGND VGND VPWR VPWR _06696_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_51_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08435_ _08470_/A _08430_/X _08431_/X _08564_/B _08434_/Y VGND VGND VPWR VPWR _08450_/C
+ sky130_fd_sc_hd__a32o_2
XFILLER_12_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08366_ _08366_/A VGND VGND VPWR VPWR _12716_/D sky130_fd_sc_hd__clkbuf_1
X_07317_ _13136_/Q _09120_/B VGND VGND VPWR VPWR _07318_/B sky130_fd_sc_hd__nor2_1
X_08297_ _08297_/A VGND VGND VPWR VPWR _13371_/D sky130_fd_sc_hd__clkbuf_1
X_07248_ _07428_/B _07243_/X _07244_/X _07246_/X _07247_/X _07327_/A VGND VGND VPWR
+ VPWR _07249_/D sky130_fd_sc_hd__mux4_2
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07179_ _07179_/A _07177_/C VGND VGND VPWR VPWR _07180_/B sky130_fd_sc_hd__or2b_1
XFILLER_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10190_ _10190_/A VGND VGND VPWR VPWR _14557_/D sky130_fd_sc_hd__inv_2
XFILLER_160_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12900_ _13274_/CLK _12900_/D hold1/X VGND VGND VPWR VPWR _12900_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13880_ _14657_/CLK hold427/X VGND VGND VPWR VPWR hold334/A sky130_fd_sc_hd__dfxtp_1
X_12831_ _14696_/CLK _12831_/D VGND VGND VPWR VPWR hold135/A sky130_fd_sc_hd__dfxtp_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _13700_/CLK _12762_/D VGND VGND VPWR VPWR hold433/A sky130_fd_sc_hd__dfxtp_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14610_/CLK _14501_/D VGND VGND VPWR VPWR _14501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11713_ _12149_/A VGND VGND VPWR VPWR _12621_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _13303_/CLK _12693_/D VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _14432_/CLK _14432_/D VGND VGND VPWR VPWR _14432_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11644_ _11644_/A VGND VGND VPWR VPWR _13997_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14363_ _14557_/CLK hold304/X VGND VGND VPWR VPWR _14363_/Q sky130_fd_sc_hd__dfxtp_1
Xinput16 data_i[23] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__buf_6
X_11575_ _11575_/A VGND VGND VPWR VPWR _13869_/D sky130_fd_sc_hd__clkbuf_1
Xinput27 hold3/X VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__buf_4
XFILLER_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13314_ _13314_/CLK hold416/X VGND VGND VPWR VPWR _13314_/Q sky130_fd_sc_hd__dfxtp_1
X_10526_ _14430_/D _13815_/Q _10526_/C VGND VGND VPWR VPWR _10531_/B sky130_fd_sc_hd__and3_1
XFILLER_156_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14294_ _14294_/CLK _14294_/D VGND VGND VPWR VPWR _14294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13245_ _14678_/CLK _13245_/D VGND VGND VPWR VPWR _13517_/D sky130_fd_sc_hd__dfxtp_1
X_10457_ hold79/A hold71/A _10461_/B _10456_/X VGND VGND VPWR VPWR _10465_/A sky130_fd_sc_hd__a31o_1
X_13176_ _13362_/CLK _13176_/D VGND VGND VPWR VPWR hold88/A sky130_fd_sc_hd__dfxtp_1
X_10388_ _10388_/A _10388_/B VGND VGND VPWR VPWR _10390_/B sky130_fd_sc_hd__xnor2_1
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12127_ _12127_/A VGND VGND VPWR VPWR _14478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12058_ _12058_/A VGND VGND VPWR VPWR _14447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11009_ _14300_/Q _14470_/Q _14226_/Q _14056_/Q _10993_/X _10995_/X VGND VGND VPWR
+ VPWR _11009_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06550_ _06550_/A _06550_/B VGND VGND VPWR VPWR _06550_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_34_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06481_ _06443_/X _06425_/X _06444_/Y _06429_/C VGND VGND VPWR VPWR _06484_/B sky130_fd_sc_hd__o22a_1
XFILLER_20_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08220_ _10310_/A _08220_/B _08220_/C VGND VGND VPWR VPWR _08226_/B sky130_fd_sc_hd__and3_1
XFILLER_21_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08151_ _08169_/A _08151_/B VGND VGND VPWR VPWR _08154_/A sky130_fd_sc_hd__or2_1
X_07102_ _07156_/A _07102_/B VGND VGND VPWR VPWR _07102_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_158_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08082_ _12977_/Q _13277_/Q _08084_/S VGND VGND VPWR VPWR _08083_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07033_ _07038_/A _07038_/B VGND VGND VPWR VPWR _07034_/B sky130_fd_sc_hd__xnor2_1
XFILLER_146_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14750__61 VGND VGND VPWR VPWR _14750__61/HI data_o[24] sky130_fd_sc_hd__conb_1
XFILLER_102_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08984_ _08984_/A _08984_/B _08984_/C VGND VGND VPWR VPWR _08985_/B sky130_fd_sc_hd__and3_1
XFILLER_103_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07935_ _13270_/Q _07955_/B VGND VGND VPWR VPWR _07944_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07866_ _07860_/A _07860_/B _07885_/A VGND VGND VPWR VPWR _07866_/X sky130_fd_sc_hd__o21ba_1
X_09605_ _13400_/Q _13598_/Q _09609_/S VGND VGND VPWR VPWR _09606_/A sky130_fd_sc_hd__mux2_2
X_06817_ _07878_/B _07878_/C _13009_/Q VGND VGND VPWR VPWR _06825_/C sky130_fd_sc_hd__a21oi_1
XFILLER_28_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07797_ _07797_/A _07797_/B VGND VGND VPWR VPWR _07797_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_25_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09536_ _13609_/Q _13610_/Q _13611_/Q _13612_/Q _09562_/B VGND VGND VPWR VPWR _09536_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_83_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06748_ _06852_/A _06746_/X _06747_/Y VGND VGND VPWR VPWR _06863_/B sky130_fd_sc_hd__o21ba_1
XFILLER_25_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09467_ _09467_/A _09467_/B VGND VGND VPWR VPWR _09468_/B sky130_fd_sc_hd__nor2_1
X_06679_ _07813_/B VGND VGND VPWR VPWR _07821_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08418_ hold467/X _13385_/Q _08418_/S VGND VGND VPWR VPWR _08419_/A sky130_fd_sc_hd__mux2_1
X_09398_ _08784_/X _09396_/Y _09397_/X _08532_/X VGND VGND VPWR VPWR _13594_/D sky130_fd_sc_hd__a31o_1
X_08349_ _08349_/A VGND VGND VPWR VPWR _12709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11360_ _13775_/Q _11359_/X _11376_/S VGND VGND VPWR VPWR _11361_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10311_ _10309_/Y _10311_/B VGND VGND VPWR VPWR _10312_/B sky130_fd_sc_hd__and2b_1
XFILLER_137_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11291_ _14697_/Q VGND VGND VPWR VPWR _11291_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13030_ _13294_/CLK _13030_/D hold1/X VGND VGND VPWR VPWR _13030_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10242_ _14370_/Q _10230_/X _10237_/A VGND VGND VPWR VPWR _10242_/X sky130_fd_sc_hd__a21o_1
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10173_ _10164_/X _10172_/X _14293_/D VGND VGND VPWR VPWR _10173_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13932_ _14179_/CLK hold350/X VGND VGND VPWR VPWR hold370/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13863_ _14075_/CLK _13863_/D VGND VGND VPWR VPWR _13863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12814_ _13635_/CLK _12814_/D VGND VGND VPWR VPWR hold406/A sky130_fd_sc_hd__dfxtp_1
X_13794_ _13945_/CLK _13794_/D VGND VGND VPWR VPWR _13794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _13702_/CLK _12745_/D VGND VGND VPWR VPWR hold183/A sky130_fd_sc_hd__dfxtp_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _13256_/CLK _12676_/D VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__dfxtp_1
X_14415_ _14424_/CLK _14415_/D VGND VGND VPWR VPWR _14415_/Q sky130_fd_sc_hd__dfxtp_1
X_11627_ _11627_/A VGND VGND VPWR VPWR _13989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14346_ _14357_/CLK hold227/X VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__dfxtp_1
X_11558_ _11558_/A VGND VGND VPWR VPWR _13861_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10509_ _10509_/A VGND VGND VPWR VPWR _10510_/B sky130_fd_sc_hd__inv_2
XFILLER_6_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14277_ _14724_/CLK _14277_/D VGND VGND VPWR VPWR _14277_/Q sky130_fd_sc_hd__dfxtp_1
X_11489_ _13831_/Q _11488_/X _11495_/S VGND VGND VPWR VPWR _11490_/A sky130_fd_sc_hd__mux2_1
X_13228_ _13605_/CLK hold514/X VGND VGND VPWR VPWR _13228_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _13552_/CLK _13159_/D _12609_/A VGND VGND VPWR VPWR _13159_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05981_ _11529_/B VGND VGND VPWR VPWR _14163_/D sky130_fd_sc_hd__inv_2
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07720_ _07720_/A VGND VGND VPWR VPWR _13660_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07651_ _07651_/A _07651_/B VGND VGND VPWR VPWR _07664_/B sky130_fd_sc_hd__xnor2_1
XFILLER_65_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06602_ _12900_/Q _06607_/D VGND VGND VPWR VPWR _06604_/A sky130_fd_sc_hd__and2_1
XFILLER_25_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07582_ _07583_/B _07583_/C _07583_/A VGND VGND VPWR VPWR _07582_/X sky130_fd_sc_hd__a21o_1
X_09321_ _13298_/Q _13536_/Q _09321_/S VGND VGND VPWR VPWR _09322_/A sky130_fd_sc_hd__mux2_1
X_06533_ _12888_/Q _06534_/B VGND VGND VPWR VPWR _06535_/A sky130_fd_sc_hd__and2_1
XFILLER_34_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09252_ _09255_/B _09252_/B VGND VGND VPWR VPWR _09252_/X sky130_fd_sc_hd__xor2_1
X_06464_ _06452_/A _06452_/B _06449_/A VGND VGND VPWR VPWR _06465_/B sky130_fd_sc_hd__o21bai_1
XFILLER_138_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08203_ _08193_/A _08193_/B _08189_/A VGND VGND VPWR VPWR _08204_/B sky130_fd_sc_hd__o21bai_1
X_09183_ _13537_/Q _09183_/B VGND VGND VPWR VPWR _09186_/A sky130_fd_sc_hd__nand2_1
X_06395_ _06469_/A _14432_/Q VGND VGND VPWR VPWR _06395_/X sky130_fd_sc_hd__and2b_1
X_08134_ _13356_/Q _08135_/B VGND VGND VPWR VPWR _08136_/A sky130_fd_sc_hd__or2_1
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08065_ _12969_/Q _13269_/Q _08073_/S VGND VGND VPWR VPWR _08066_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07016_ _07040_/A _07119_/A _07063_/B _07031_/A VGND VGND VPWR VPWR _07019_/A sky130_fd_sc_hd__a22oi_1
XFILLER_161_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08967_ _08967_/A _08965_/C VGND VGND VPWR VPWR _08968_/B sky130_fd_sc_hd__or2b_1
XFILLER_124_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07918_ _07898_/A _07904_/A _07905_/A VGND VGND VPWR VPWR _07918_/Y sky130_fd_sc_hd__o21bai_1
X_08898_ _13428_/Q _13429_/Q _08929_/C _13520_/D VGND VGND VPWR VPWR _08899_/B sky130_fd_sc_hd__and4_1
XFILLER_84_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07849_ _07858_/C _07842_/B _07848_/Y VGND VGND VPWR VPWR _07850_/B sky130_fd_sc_hd__o21ai_1
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10860_ _10860_/A VGND VGND VPWR VPWR _13189_/D sky130_fd_sc_hd__clkbuf_1
X_09519_ _09519_/A _09519_/B VGND VGND VPWR VPWR _09534_/B sky130_fd_sc_hd__nand2_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10791_ _10791_/A VGND VGND VPWR VPWR _13058_/D sky130_fd_sc_hd__clkbuf_1
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _11307_/X _14711_/Q _12532_/S VGND VGND VPWR VPWR _12531_/A sky130_fd_sc_hd__mux2_1
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12461_ _14662_/Q _14519_/Q _12461_/S VGND VGND VPWR VPWR _12462_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14200_ _14210_/CLK _14200_/D VGND VGND VPWR VPWR _14200_/Q sky130_fd_sc_hd__dfxtp_1
X_11412_ _13729_/Q _11416_/B VGND VGND VPWR VPWR _11413_/A sky130_fd_sc_hd__and2_1
XFILLER_149_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12392_ _14618_/Q _12022_/X _12394_/S VGND VGND VPWR VPWR _12393_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14131_ _14716_/CLK hold412/X VGND VGND VPWR VPWR hold241/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11343_ _12007_/A VGND VGND VPWR VPWR _11343_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14062_ _14543_/CLK _14062_/D VGND VGND VPWR VPWR _14062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11274_ _14728_/Q VGND VGND VPWR VPWR _11274_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13013_ _13303_/CLK _13013_/D repeater59/X VGND VGND VPWR VPWR _13013_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10225_ _10225_/A VGND VGND VPWR VPWR _14400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10156_ _14284_/D _10155_/X _14294_/D VGND VGND VPWR VPWR _10157_/A sky130_fd_sc_hd__mux2_1
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_10087_ _10082_/X _10086_/X _14048_/D VGND VGND VPWR VPWR _10088_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13915_ _14047_/CLK hold160/X VGND VGND VPWR VPWR hold197/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13846_ _14042_/CLK hold156/X VGND VGND VPWR VPWR hold97/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13777_ _14725_/CLK _13777_/D VGND VGND VPWR VPWR _13777_/Q sky130_fd_sc_hd__dfxtp_1
X_10989_ _11037_/A _10989_/B VGND VGND VPWR VPWR _10989_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12728_ _13372_/CLK _12728_/D VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12659_ _14737_/CLK hold403/X _12609_/A VGND VGND VPWR VPWR hold488/A sky130_fd_sc_hd__dfrtp_1
XFILLER_129_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06180_ _13847_/Q _13848_/Q _13849_/Q _13850_/Q VGND VGND VPWR VPWR _06180_/X sky130_fd_sc_hd__or4_1
XFILLER_116_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14329_ _14696_/CLK hold398/X VGND VGND VPWR VPWR hold364/A sky130_fd_sc_hd__dfxtp_1
Xhold405 hold405/A VGND VGND VPWR VPWR hold405/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold416 hold416/A VGND VGND VPWR VPWR hold416/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold427 hold427/A VGND VGND VPWR VPWR hold427/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold438 hold438/A VGND VGND VPWR VPWR hold438/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold449 hold449/A VGND VGND VPWR VPWR hold449/X sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _13689_/Q _09870_/B _09873_/D VGND VGND VPWR VPWR _09872_/A sky130_fd_sc_hd__and3_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _08826_/A _08826_/B VGND VGND VPWR VPWR _08822_/B sky130_fd_sc_hd__xnor2_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08752_ _09576_/B VGND VGND VPWR VPWR _09581_/B sky130_fd_sc_hd__buf_2
XFILLER_97_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05964_ _14075_/D _13630_/Q _05957_/X _05959_/X _05963_/Y VGND VGND VPWR VPWR _05979_/A
+ sky130_fd_sc_hd__a41o_1
XFILLER_39_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07703_ _07703_/A _07703_/B VGND VGND VPWR VPWR _07705_/C sky130_fd_sc_hd__xnor2_1
XFILLER_38_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08683_ _09506_/A VGND VGND VPWR VPWR _09493_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07634_ _07635_/A _07635_/B VGND VGND VPWR VPWR _07659_/B sky130_fd_sc_hd__and2_1
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07565_ _13159_/Q _09271_/B VGND VGND VPWR VPWR _07566_/B sky130_fd_sc_hd__nor2_1
XFILLER_22_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09304_ _13290_/Q _13528_/Q _09310_/S VGND VGND VPWR VPWR _09305_/A sky130_fd_sc_hd__mux2_1
X_06516_ _06516_/A VGND VGND VPWR VPWR _06519_/A sky130_fd_sc_hd__inv_2
X_07496_ _13150_/Q _07513_/B VGND VGND VPWR VPWR _07504_/D sky130_fd_sc_hd__xnor2_1
XFILLER_10_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09235_ _09230_/A _09228_/X _09241_/A _09229_/A VGND VGND VPWR VPWR _09235_/X sky130_fd_sc_hd__a211o_1
X_06447_ _12880_/Q _06448_/B VGND VGND VPWR VPWR _06449_/A sky130_fd_sc_hd__and2_1
XFILLER_10_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09166_ _09158_/X _09160_/X _09162_/X _09165_/Y VGND VGND VPWR VPWR _09173_/B sky130_fd_sc_hd__a31o_1
X_06378_ _06429_/A VGND VGND VPWR VPWR _06446_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08117_ _13477_/Q _14011_/Q _14009_/Q _14007_/Q _08142_/A _08143_/A VGND VGND VPWR
+ VPWR _08220_/C sky130_fd_sc_hd__mux4_2
X_09097_ _07570_/X _09095_/X _09096_/Y _07279_/X VGND VGND VPWR VPWR _13525_/D sky130_fd_sc_hd__a31o_1
XFILLER_134_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08048_ _08048_/A VGND VGND VPWR VPWR _12685_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10010_ _13909_/Q VGND VGND VPWR VPWR _10052_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_131_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09999_ _09994_/X _11270_/B _10635_/B VGND VGND VPWR VPWR _10000_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11961_ _11961_/A VGND VGND VPWR VPWR _14297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10912_ _11186_/A VGND VGND VPWR VPWR _12586_/A sky130_fd_sc_hd__clkbuf_4
X_13700_ _13700_/CLK _13700_/D VGND VGND VPWR VPWR _13700_/Q sky130_fd_sc_hd__dfxtp_2
X_14680_ _14680_/CLK _14680_/D VGND VGND VPWR VPWR hold442/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11892_ _14243_/Q _11519_/X _11894_/S VGND VGND VPWR VPWR _11893_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13631_ _13855_/CLK hold466/X VGND VGND VPWR VPWR _13631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10843_ _10876_/A VGND VGND VPWR VPWR _10852_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_71_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13562_ _13562_/CLK hold192/X VGND VGND VPWR VPWR _13562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10774_ _10774_/A VGND VGND VPWR VPWR _13050_/D sky130_fd_sc_hd__clkbuf_1
X_12513_ _11272_/X _14703_/Q _12521_/S VGND VGND VPWR VPWR _12514_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13493_ _13704_/CLK hold259/X VGND VGND VPWR VPWR _13493_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_160_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _14697_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_12_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12444_ _14654_/Q _14700_/Q _12450_/S VGND VGND VPWR VPWR _12445_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12375_ _14610_/Q _11997_/X _12375_/S VGND VGND VPWR VPWR _12376_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14114_ _14693_/CLK hold37/X VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__dfxtp_1
X_11326_ _14519_/Q VGND VGND VPWR VPWR _11326_/X sky130_fd_sc_hd__buf_2
XFILLER_153_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14045_ _14050_/CLK _14045_/D VGND VGND VPWR VPWR _14045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11257_ _11257_/A _10960_/A VGND VGND VPWR VPWR _11257_/X sky130_fd_sc_hd__or2b_1
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10208_ _06226_/X _06325_/X _10208_/S VGND VGND VPWR VPWR _10209_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11188_ _14613_/Q _14575_/Q _14506_/Q _14458_/Q _11186_/X _11187_/X VGND VGND VPWR
+ VPWR _11189_/A sky130_fd_sc_hd__mux4_1
XFILLER_95_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10139_ _10139_/A _14160_/Q VGND VGND VPWR VPWR _10149_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13829_ _14713_/CLK _13829_/D VGND VGND VPWR VPWR _13829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07350_ _07350_/A _07375_/B VGND VGND VPWR VPWR _07364_/A sky130_fd_sc_hd__nand2_2
X_06301_ _13871_/Q _13855_/Q _06309_/S VGND VGND VPWR VPWR _06302_/A sky130_fd_sc_hd__mux2_1
X_07281_ _13169_/Q _13664_/Q _13666_/Q _13662_/Q _07247_/X _07267_/S VGND VGND VPWR
+ VPWR _07400_/B sky130_fd_sc_hd__mux4_2
Xclkbuf_leaf_151_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _14543_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09020_ _09655_/S VGND VGND VPWR VPWR _09029_/S sky130_fd_sc_hd__clkbuf_2
X_06232_ _14087_/Q _06245_/B VGND VGND VPWR VPWR _06233_/A sky130_fd_sc_hd__and2_1
XFILLER_164_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06163_ _06163_/A VGND VGND VPWR VPWR _14169_/D sky130_fd_sc_hd__clkbuf_1
Xhold202 hold202/A VGND VGND VPWR VPWR hold202/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_145_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold213 hold213/A VGND VGND VPWR VPWR hold213/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold224 hold224/A VGND VGND VPWR VPWR hold224/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold235 hold235/A VGND VGND VPWR VPWR hold235/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06094_ _06105_/B VGND VGND VPWR VPWR _11593_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold246 hold246/A VGND VGND VPWR VPWR hold246/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold257 hold257/A VGND VGND VPWR VPWR hold257/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold268 hold268/A VGND VGND VPWR VPWR hold268/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold279 hold279/A VGND VGND VPWR VPWR hold279/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09922_ _13486_/Q _13675_/Q _09924_/S VGND VGND VPWR VPWR _09923_/A sky130_fd_sc_hd__mux2_1
X_09853_ _09851_/X _09894_/A _09853_/C VGND VGND VPWR VPWR _09854_/A sky130_fd_sc_hd__and3b_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08804_ _08828_/A _08907_/A _08851_/B _08819_/A VGND VGND VPWR VPWR _08807_/A sky130_fd_sc_hd__a22oi_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _09855_/A VGND VGND VPWR VPWR _09894_/A sky130_fd_sc_hd__buf_2
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06996_ _06996_/A _06996_/B _06990_/Y _06991_/X VGND VGND VPWR VPWR _07001_/C sky130_fd_sc_hd__or4bb_1
XFILLER_105_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ _09506_/A VGND VGND VPWR VPWR _08735_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05947_ _13875_/Q _13876_/Q _13877_/Q VGND VGND VPWR VPWR _05950_/A sky130_fd_sc_hd__and3_1
XFILLER_73_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ _08617_/X _08663_/X _08664_/Y _08665_/X VGND VGND VPWR VPWR _13450_/D sky130_fd_sc_hd__a31o_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07617_ _07602_/Y _07616_/Y _11266_/A VGND VGND VPWR VPWR _07618_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08597_ _08607_/A _08605_/A VGND VGND VPWR VPWR _08602_/A sky130_fd_sc_hd__xnor2_1
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07548_ _07548_/A _07548_/B VGND VGND VPWR VPWR _07553_/C sky130_fd_sc_hd__nand2_1
XFILLER_139_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_142_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _14209_/CLK sky130_fd_sc_hd__clkbuf_16
X_07479_ _09207_/B VGND VGND VPWR VPWR _09228_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09218_ _13543_/Q _09237_/B VGND VGND VPWR VPWR _09219_/B sky130_fd_sc_hd__nor2_1
XFILLER_139_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10490_ _10490_/A _10490_/B _10490_/C VGND VGND VPWR VPWR _10491_/B sky130_fd_sc_hd__or3_1
XFILLER_154_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09149_ _09159_/A _09149_/B VGND VGND VPWR VPWR _09149_/Y sky130_fd_sc_hd__nand2_1
X_12160_ _12160_/A VGND VGND VPWR VPWR _14492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11111_ _14025_/Q _13991_/Q _13831_/Q _14543_/Q _11081_/X _11082_/X VGND VGND VPWR
+ VPWR _11112_/A sky130_fd_sc_hd__mux4_1
XFILLER_162_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12091_ _11370_/X _14463_/Q _12093_/S VGND VGND VPWR VPWR _12092_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11042_ _10991_/X _11039_/X _11041_/X _11015_/X VGND VGND VPWR VPWR _11042_/X sky130_fd_sc_hd__o211a_1
XFILLER_39_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12993_ _14633_/CLK _13815_/Q VGND VGND VPWR VPWR _13115_/D sky130_fd_sc_hd__dfxtp_2
X_14732_ _14732_/CLK _14732_/D VGND VGND VPWR VPWR _14732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11944_ _14278_/Q _11516_/X _11948_/S VGND VGND VPWR VPWR _11945_/A sky130_fd_sc_hd__mux2_1
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11875_ _14235_/Q _11494_/X _11875_/S VGND VGND VPWR VPWR _11876_/A sky130_fd_sc_hd__mux2_1
X_14663_ _14667_/CLK _14663_/D VGND VGND VPWR VPWR _14663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13614_ _13635_/CLK _13614_/D repeater57/X VGND VGND VPWR VPWR _13614_/Q sky130_fd_sc_hd__dfrtp_2
X_10826_ _10826_/A VGND VGND VPWR VPWR _13174_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14594_ _14643_/CLK _14594_/D VGND VGND VPWR VPWR _14594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13545_ _13587_/CLK _13545_/D _12609_/A VGND VGND VPWR VPWR _13545_/Q sky130_fd_sc_hd__dfrtp_2
X_10757_ _13001_/Q _10820_/A VGND VGND VPWR VPWR _10758_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_133_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _14201_/CLK sky130_fd_sc_hd__clkbuf_16
X_13476_ _13476_/CLK _13476_/D VGND VGND VPWR VPWR _13476_/Q sky130_fd_sc_hd__dfxtp_1
X_10688_ _10688_/A VGND VGND VPWR VPWR _12923_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12427_ _12427_/A VGND VGND VPWR VPWR _14646_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12358_ _14602_/Q _11972_/X _12364_/S VGND VGND VPWR VPWR _12359_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11309_ _11309_/A VGND VGND VPWR VPWR _13763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12289_ _14561_/Q _11962_/X _12291_/S VGND VGND VPWR VPWR _12290_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14028_ _14720_/CLK _14028_/D VGND VGND VPWR VPWR _14028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06850_ _06665_/X _06847_/Y _06848_/X _06849_/X VGND VGND VPWR VPWR _13011_/D sky130_fd_sc_hd__a31o_1
XFILLER_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06781_ _13006_/Q _06781_/B VGND VGND VPWR VPWR _06794_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08520_ _08535_/A _08520_/B _08520_/C VGND VGND VPWR VPWR _08552_/A sky130_fd_sc_hd__and3_1
XFILLER_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08451_ _08490_/A VGND VGND VPWR VPWR _09367_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07402_ _07461_/C VGND VGND VPWR VPWR _09153_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_08382_ _13088_/Q _13369_/Q _08384_/S VGND VGND VPWR VPWR _08383_/A sky130_fd_sc_hd__mux2_1
X_07333_ _07387_/A _07333_/B VGND VGND VPWR VPWR _07333_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_124_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _13811_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07264_ _07299_/S VGND VGND VPWR VPWR _07267_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09003_ _09003_/A _09003_/B VGND VGND VPWR VPWR _09003_/Y sky130_fd_sc_hd__xnor2_1
X_06215_ _14379_/Q _06324_/A _06215_/C _06215_/D VGND VGND VPWR VPWR _06216_/B sky130_fd_sc_hd__or4_1
XFILLER_118_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07195_ _07196_/A _07196_/B _07196_/C VGND VGND VPWR VPWR _07197_/A sky130_fd_sc_hd__a21oi_1
XFILLER_145_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06146_ _06146_/A _06146_/B VGND VGND VPWR VPWR _06146_/Y sky130_fd_sc_hd__nor2_1
XFILLER_160_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06077_ _06259_/A _06259_/B _06076_/Y VGND VGND VPWR VPWR _06257_/S sky130_fd_sc_hd__a21oi_1
XFILLER_132_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09905_ _13478_/Q _13667_/Q _09913_/S VGND VGND VPWR VPWR _09906_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09836_ _09836_/A _09836_/B _14440_/Q _09836_/D VGND VGND VPWR VPWR _09838_/B sky130_fd_sc_hd__and4_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06979_ _06981_/B _06979_/B VGND VGND VPWR VPWR _06979_/Y sky130_fd_sc_hd__xnor2_1
X_09767_ _09767_/A _13703_/Q VGND VGND VPWR VPWR _09809_/C sky130_fd_sc_hd__nor2_2
XFILLER_55_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _08741_/A _08718_/B VGND VGND VPWR VPWR _08718_/X sky130_fd_sc_hd__xor2_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _09695_/B _09697_/Y _09883_/B VGND VGND VPWR VPWR _09699_/A sky130_fd_sc_hd__mux2_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _13449_/Q _09464_/B VGND VGND VPWR VPWR _08664_/A sky130_fd_sc_hd__nand2_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11660_ _11660_/A VGND VGND VPWR VPWR _14013_/D sky130_fd_sc_hd__clkbuf_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10611_ _14044_/Q _14043_/Q VGND VGND VPWR VPWR _10611_/X sky130_fd_sc_hd__or2_1
XFILLER_23_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11591_ _14075_/D _11591_/B VGND VGND VPWR VPWR _11592_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_115_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _13619_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13330_ _14610_/CLK _13330_/D VGND VGND VPWR VPWR _13330_/Q sky130_fd_sc_hd__dfxtp_2
X_10542_ _10542_/A _10542_/B VGND VGND VPWR VPWR _14435_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13261_ _13263_/CLK _13261_/D hold1/X VGND VGND VPWR VPWR _13261_/Q sky130_fd_sc_hd__dfrtp_1
X_10473_ _10495_/A _10485_/A _10485_/B hold186/A VGND VGND VPWR VPWR _10474_/A sky130_fd_sc_hd__a22o_1
X_12212_ _14122_/Q _12215_/C VGND VGND VPWR VPWR _12214_/A sky130_fd_sc_hd__and2_1
XFILLER_124_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13192_ _13606_/CLK _13192_/D VGND VGND VPWR VPWR hold509/A sky130_fd_sc_hd__dfxtp_1
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12143_ _14486_/Q _12019_/X _12147_/S VGND VGND VPWR VPWR _12144_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12074_ _11326_/X _14455_/Q _12074_/S VGND VGND VPWR VPWR _12075_/A sky130_fd_sc_hd__mux2_1
X_11025_ _11017_/X _11019_/Y _11023_/Y _11024_/X VGND VGND VPWR VPWR _11026_/B sky130_fd_sc_hd__a211o_1
XFILLER_37_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12976_ _13280_/CLK hold255/X VGND VGND VPWR VPWR _12976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14715_ _14717_/CLK _14715_/D VGND VGND VPWR VPWR _14715_/Q sky130_fd_sc_hd__dfxtp_1
X_11927_ _14270_/Q _11491_/X _11929_/S VGND VGND VPWR VPWR _11928_/A sky130_fd_sc_hd__mux2_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14646_ _14679_/CLK _14646_/D VGND VGND VPWR VPWR _14646_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11858_ _14227_/Q _11469_/X _11864_/S VGND VGND VPWR VPWR _11859_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_19 input26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10809_ _10809_/A VGND VGND VPWR VPWR _13066_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_106_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _13598_/CLK sky130_fd_sc_hd__clkbuf_16
X_14577_ _14579_/CLK _14577_/D VGND VGND VPWR VPWR _14577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11789_ _13566_/Q _11795_/B VGND VGND VPWR VPWR _11790_/A sky130_fd_sc_hd__and2_1
XFILLER_159_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13528_ _13528_/CLK _13528_/D _12609_/A VGND VGND VPWR VPWR _13528_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13459_ _13626_/CLK _13459_/D repeater57/X VGND VGND VPWR VPWR _13459_/Q sky130_fd_sc_hd__dfrtp_2
X_06000_ _13569_/Q _13570_/Q _13571_/Q _13576_/Q VGND VGND VPWR VPWR _06001_/D sky130_fd_sc_hd__or4_1
XFILLER_115_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07951_ _07925_/A _07973_/A _07975_/A VGND VGND VPWR VPWR _07953_/B sky130_fd_sc_hd__o21ba_1
XFILLER_141_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06902_ _07962_/B VGND VGND VPWR VPWR _07963_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_141_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07882_ _07811_/X _07880_/X _07881_/Y _06821_/X VGND VGND VPWR VPWR _13263_/D sky130_fd_sc_hd__a31o_1
XFILLER_95_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09621_ _09621_/A VGND VGND VPWR VPWR _12824_/D sky130_fd_sc_hd__clkbuf_1
X_06833_ _13010_/Q _07889_/B VGND VGND VPWR VPWR _06834_/B sky130_fd_sc_hd__or2_1
XFILLER_37_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09552_ _09553_/B _09553_/C _09559_/A VGND VGND VPWR VPWR _09556_/B sky130_fd_sc_hd__a21o_1
XFILLER_71_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06764_ _07861_/S VGND VGND VPWR VPWR _07843_/S sky130_fd_sc_hd__buf_2
XFILLER_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08503_ _08503_/A VGND VGND VPWR VPWR _13438_/D sky130_fd_sc_hd__clkbuf_1
X_09483_ _13605_/Q _09518_/B VGND VGND VPWR VPWR _09484_/B sky130_fd_sc_hd__or2_1
X_06695_ _13001_/Q _06695_/B VGND VGND VPWR VPWR _06712_/A sky130_fd_sc_hd__nor2_1
XFILLER_51_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08434_ _13471_/Q _13476_/Q VGND VGND VPWR VPWR _08434_/Y sky130_fd_sc_hd__nor2_2
XFILLER_12_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08365_ _13080_/Q _13361_/Q _08373_/S VGND VGND VPWR VPWR _08366_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07316_ _07316_/A VGND VGND VPWR VPWR _07318_/A sky130_fd_sc_hd__clkinv_2
X_08296_ _08294_/X _08296_/B _08296_/C VGND VGND VPWR VPWR _08297_/A sky130_fd_sc_hd__and3b_1
XFILLER_164_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07247_ _13171_/Q VGND VGND VPWR VPWR _07247_/X sky130_fd_sc_hd__buf_2
Xclkbuf_4_2_0_clk clkbuf_4_3_0_clk/A VGND VGND VPWR VPWR clkbuf_4_2_0_clk/X sky130_fd_sc_hd__clkbuf_2
X_07178_ _07178_/A _07178_/B VGND VGND VPWR VPWR _07179_/A sky130_fd_sc_hd__nor2_1
X_06129_ _06129_/A VGND VGND VPWR VPWR _14150_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09819_ _09836_/A _09819_/B _09836_/D VGND VGND VPWR VPWR _09821_/B sky130_fd_sc_hd__and3_1
XFILLER_143_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12830_ _13653_/CLK _12830_/D VGND VGND VPWR VPWR hold92/A sky130_fd_sc_hd__dfxtp_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _13602_/CLK _12761_/D VGND VGND VPWR VPWR hold89/A sky130_fd_sc_hd__dfxtp_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _14602_/CLK _14500_/D VGND VGND VPWR VPWR _14500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _14736_/Q _11712_/B _12564_/A VGND VGND VPWR VPWR _12041_/C sky130_fd_sc_hd__and3_2
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _13304_/CLK _12692_/D VGND VGND VPWR VPWR hold111/A sky130_fd_sc_hd__dfxtp_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _13997_/Q _11507_/X _11645_/S VGND VGND VPWR VPWR _11644_/A sky130_fd_sc_hd__mux2_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14431_ _14435_/CLK _14431_/D VGND VGND VPWR VPWR _14431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11574_ _13645_/Q _11574_/B VGND VGND VPWR VPWR _11575_/A sky130_fd_sc_hd__and2_1
X_14362_ _14425_/CLK _14362_/D VGND VGND VPWR VPWR _14362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput17 data_i[2] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__buf_6
Xinput28 rtr_i VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__buf_12
XFILLER_128_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10525_ _10525_/A _10525_/B VGND VGND VPWR VPWR _14434_/D sky130_fd_sc_hd__xor2_1
X_13313_ _14275_/CLK hold76/X VGND VGND VPWR VPWR _13313_/Q sky130_fd_sc_hd__dfxtp_1
X_14293_ _14294_/CLK _14293_/D VGND VGND VPWR VPWR _14293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13244_ _14687_/CLK _13244_/D VGND VGND VPWR VPWR _13516_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10456_ hold46/A hold62/A _10456_/C VGND VGND VPWR VPWR _10456_/X sky130_fd_sc_hd__and3_1
XFILLER_124_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13175_ _13362_/CLK _13175_/D VGND VGND VPWR VPWR hold65/A sky130_fd_sc_hd__dfxtp_1
X_10387_ _10382_/X _10387_/B VGND VGND VPWR VPWR _10388_/B sky130_fd_sc_hd__and2b_1
XFILLER_124_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12126_ _14478_/Q _11994_/X _12128_/S VGND VGND VPWR VPWR _12127_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12057_ _11301_/X _14447_/Q _12063_/S VGND VGND VPWR VPWR _12058_/A sky130_fd_sc_hd__mux2_1
X_11008_ _12645_/B VGND VGND VPWR VPWR _11008_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12959_ _13263_/CLK hold91/X VGND VGND VPWR VPWR _12959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06480_ _06480_/A VGND VGND VPWR VPWR _12882_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14629_ _14645_/CLK hold486/X VGND VGND VPWR VPWR _14629_/Q sky130_fd_sc_hd__dfxtp_1
X_08150_ _13357_/Q _08150_/B VGND VGND VPWR VPWR _08151_/B sky130_fd_sc_hd__and2_1
XFILLER_158_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07101_ _07101_/A _07101_/B VGND VGND VPWR VPWR _07102_/B sky130_fd_sc_hd__xnor2_1
XFILLER_119_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08081_ _08081_/A VGND VGND VPWR VPWR _12700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07032_ _07032_/A _07032_/B VGND VGND VPWR VPWR _07038_/B sky130_fd_sc_hd__xnor2_1
XFILLER_162_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08983_ _08984_/A _08984_/B _08984_/C VGND VGND VPWR VPWR _08985_/A sky130_fd_sc_hd__a21oi_1
XFILLER_142_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07934_ _07934_/A _07930_/B VGND VGND VPWR VPWR _07939_/B sky130_fd_sc_hd__or2b_1
XFILLER_68_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07865_ _07885_/D VGND VGND VPWR VPWR _07892_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09604_ _09604_/A VGND VGND VPWR VPWR _12816_/D sky130_fd_sc_hd__clkbuf_1
X_06816_ _13009_/Q _07878_/B _07878_/C VGND VGND VPWR VPWR _06825_/B sky130_fd_sc_hd__and3_1
X_07796_ _07796_/A _07796_/B VGND VGND VPWR VPWR _07797_/B sky130_fd_sc_hd__xnor2_1
XFILLER_44_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09535_ _09535_/A _09535_/B VGND VGND VPWR VPWR _09535_/X sky130_fd_sc_hd__or2_1
X_06747_ _06783_/S _13036_/Q VGND VGND VPWR VPWR _06747_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09466_ _09466_/A _09466_/B VGND VGND VPWR VPWR _09467_/B sky130_fd_sc_hd__nor2_1
X_06678_ _13000_/Q _07813_/B VGND VGND VPWR VPWR _06681_/B sky130_fd_sc_hd__nor2_1
X_08417_ _08417_/A VGND VGND VPWR VPWR _12739_/D sky130_fd_sc_hd__clkbuf_1
X_09397_ _09396_/A _09419_/A _09419_/B VGND VGND VPWR VPWR _09397_/X sky130_fd_sc_hd__a21o_1
XFILLER_11_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08348_ _13073_/Q _13354_/Q _10891_/B VGND VGND VPWR VPWR _08349_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08279_ _10304_/A _10306_/A _13477_/Q _08279_/D VGND VGND VPWR VPWR _08281_/B sky130_fd_sc_hd__and4_1
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10310_ _10310_/A _13513_/D VGND VGND VPWR VPWR _10311_/B sky130_fd_sc_hd__nand2_1
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11290_ _11290_/A VGND VGND VPWR VPWR _13757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10241_ _14366_/Q _10230_/X _10237_/A VGND VGND VPWR VPWR _14523_/D sky130_fd_sc_hd__a21o_1
XFILLER_105_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10172_ _10103_/A _10150_/X _10159_/X VGND VGND VPWR VPWR _10172_/X sky130_fd_sc_hd__a21o_1
XFILLER_79_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13931_ _14179_/CLK _13931_/D VGND VGND VPWR VPWR hold350/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13862_ _14075_/CLK _13862_/D VGND VGND VPWR VPWR _13862_/Q sky130_fd_sc_hd__dfxtp_1
X_12813_ _13635_/CLK _12813_/D VGND VGND VPWR VPWR hold381/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13793_ _13799_/CLK _13793_/D VGND VGND VPWR VPWR _13793_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _13702_/CLK _12744_/D VGND VGND VPWR VPWR hold185/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _13525_/CLK _12675_/D VGND VGND VPWR VPWR hold233/A sky130_fd_sc_hd__dfxtp_1
X_14414_ _14424_/CLK _14414_/D VGND VGND VPWR VPWR hold354/A sky130_fd_sc_hd__dfxtp_1
X_11626_ _13989_/Q _11481_/X _11634_/S VGND VGND VPWR VPWR _11627_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14345_ _14697_/CLK hold490/X VGND VGND VPWR VPWR hold113/A sky130_fd_sc_hd__dfxtp_1
X_11557_ _13637_/Q _11563_/B VGND VGND VPWR VPWR _11558_/A sky130_fd_sc_hd__and2_1
XFILLER_116_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10508_ _12989_/D VGND VGND VPWR VPWR _10509_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11488_ _14517_/Q VGND VGND VPWR VPWR _11488_/X sky130_fd_sc_hd__clkbuf_2
X_14276_ _14667_/CLK _14276_/D VGND VGND VPWR VPWR _14276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13227_ _13605_/CLK hold521/X VGND VGND VPWR VPWR _13227_/Q sky130_fd_sc_hd__dfxtp_1
X_10439_ _10439_/A _14004_/D VGND VGND VPWR VPWR _10439_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _14530_/CLK _13158_/D _12609_/A VGND VGND VPWR VPWR _13158_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _14470_/Q _11968_/X _12117_/S VGND VGND VPWR VPWR _12110_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05980_ _11576_/A VGND VGND VPWR VPWR _11529_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13089_ _13558_/CLK hold108/X VGND VGND VPWR VPWR _13089_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07650_ _14702_/Q _13114_/Q VGND VGND VPWR VPWR _07651_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06601_ _06607_/D _06601_/B VGND VGND VPWR VPWR _12899_/D sky130_fd_sc_hd__nor2_1
XFILLER_65_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07581_ _07581_/A _07581_/B VGND VGND VPWR VPWR _07583_/A sky130_fd_sc_hd__or2_1
X_09320_ _09320_/A VGND VGND VPWR VPWR _12787_/D sky130_fd_sc_hd__clkbuf_1
X_06532_ _06543_/A _06532_/B _06554_/C VGND VGND VPWR VPWR _06534_/B sky130_fd_sc_hd__and3_1
XFILLER_22_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09251_ _13547_/Q _09289_/B _09256_/A _09255_/A VGND VGND VPWR VPWR _09252_/B sky130_fd_sc_hd__a22o_1
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06463_ _06463_/A _06462_/X VGND VGND VPWR VPWR _06465_/A sky130_fd_sc_hd__or2b_1
XFILLER_22_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08202_ _08202_/A _08202_/B VGND VGND VPWR VPWR _08204_/A sky130_fd_sc_hd__or2_1
X_09182_ _09182_/A VGND VGND VPWR VPWR _09182_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06394_ _13106_/D VGND VGND VPWR VPWR _06469_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08133_ _08123_/A _08121_/X _08122_/A VGND VGND VPWR VPWR _08137_/A sky130_fd_sc_hd__a21o_1
XFILLER_162_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08064_ _08097_/A VGND VGND VPWR VPWR _08073_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_135_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07015_ hold515/A VGND VGND VPWR VPWR _07063_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08966_ _08966_/A _08966_/B VGND VGND VPWR VPWR _08967_/A sky130_fd_sc_hd__nor2_1
XFILLER_57_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07917_ _07917_/A _07917_/B VGND VGND VPWR VPWR _07917_/Y sky130_fd_sc_hd__nand2_1
X_08897_ _13429_/Q _08929_/C _08951_/B _13428_/Q VGND VGND VPWR VPWR _08899_/A sky130_fd_sc_hd__a22oi_1
XFILLER_29_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_95_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _13721_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07848_ _13258_/Q _07856_/B VGND VGND VPWR VPWR _07848_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07779_ _07779_/A _07779_/B VGND VGND VPWR VPWR _07780_/B sky130_fd_sc_hd__or2_1
XFILLER_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09518_ _13610_/Q _09518_/B VGND VGND VPWR VPWR _09519_/B sky130_fd_sc_hd__or2_1
X_10790_ _13016_/Q _10790_/B VGND VGND VPWR VPWR _10791_/A sky130_fd_sc_hd__and2_1
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09449_ _09420_/A _09420_/B _09420_/C _09420_/D _09448_/Y VGND VGND VPWR VPWR _09449_/Y
+ sky130_fd_sc_hd__o41ai_2
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12460_ _12460_/A VGND VGND VPWR VPWR _14661_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11411_ _11411_/A VGND VGND VPWR VPWR _13797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12391_ _12391_/A VGND VGND VPWR VPWR _14617_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11342_ _11351_/C _11353_/B _11342_/C VGND VGND VPWR VPWR _12007_/A sky130_fd_sc_hd__and3b_4
X_14130_ _14159_/CLK hold292/X VGND VGND VPWR VPWR hold237/A sky130_fd_sc_hd__dfxtp_1
XFILLER_137_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11273_ _14735_/Q VGND VGND VPWR VPWR _11712_/B sky130_fd_sc_hd__clkbuf_2
X_14061_ _14543_/CLK _14061_/D VGND VGND VPWR VPWR _14061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10224_ _14101_/Q _14085_/Q _10224_/S VGND VGND VPWR VPWR _10225_/A sky130_fd_sc_hd__mux2_1
X_13012_ _13303_/CLK _13012_/D repeater59/X VGND VGND VPWR VPWR _13012_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10155_ _14153_/Q _10143_/X _10150_/A VGND VGND VPWR VPWR _10155_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10086_ _10077_/X _10085_/X _14049_/D VGND VGND VPWR VPWR _10086_/X sky130_fd_sc_hd__mux2_1
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_87_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_86_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _14256_/CLK sky130_fd_sc_hd__clkbuf_16
X_13914_ _14047_/CLK hold197/X VGND VGND VPWR VPWR _13914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13845_ _14196_/CLK hold97/X VGND VGND VPWR VPWR hold146/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13776_ _14724_/CLK _13776_/D VGND VGND VPWR VPWR _13776_/Q sky130_fd_sc_hd__dfxtp_1
X_10988_ _10932_/X _10985_/Y _10987_/Y _10946_/X VGND VGND VPWR VPWR _10989_/B sky130_fd_sc_hd__a211o_1
XFILLER_16_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12727_ _13372_/CLK _12727_/D VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12658_ _14555_/CLK hold510/X _12609_/A VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__dfrtp_1
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11609_ _11609_/A VGND VGND VPWR VPWR _13981_/D sky130_fd_sc_hd__clkbuf_1
X_12589_ _14749_/Q _14734_/Q VGND VGND VPWR VPWR _12591_/C sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_10_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _13283_/CLK sky130_fd_sc_hd__clkbuf_16
X_14328_ _14696_/CLK hold364/X VGND VGND VPWR VPWR hold140/A sky130_fd_sc_hd__dfxtp_1
XFILLER_117_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold406 hold406/A VGND VGND VPWR VPWR hold406/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_128_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold417 hold417/A VGND VGND VPWR VPWR hold417/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold428 hold428/A VGND VGND VPWR VPWR hold428/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold439 hold439/A VGND VGND VPWR VPWR hold439/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14259_ _14707_/CLK _14259_/D VGND VGND VPWR VPWR _14259_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _08820_/A _08820_/B VGND VGND VPWR VPWR _08826_/B sky130_fd_sc_hd__xnor2_1
XFILLER_98_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05963_ _14075_/D _13630_/Q _05963_/C _05963_/D VGND VGND VPWR VPWR _05963_/Y sky130_fd_sc_hd__nor4_1
X_08751_ _13460_/Q _09542_/B VGND VGND VPWR VPWR _08757_/B sky130_fd_sc_hd__xor2_1
XFILLER_112_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _13657_/CLK sky130_fd_sc_hd__clkbuf_16
X_07702_ _07702_/A _07732_/A VGND VGND VPWR VPWR _07703_/B sky130_fd_sc_hd__nor2_1
X_08682_ _08682_/A _08787_/B VGND VGND VPWR VPWR _09506_/A sky130_fd_sc_hd__and2_1
X_07633_ _07640_/B _07633_/B VGND VGND VPWR VPWR _07635_/B sky130_fd_sc_hd__xnor2_1
XFILLER_19_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07564_ _13159_/Q _09271_/B VGND VGND VPWR VPWR _07566_/A sky130_fd_sc_hd__and2_1
XFILLER_110_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09303_ _09303_/A VGND VGND VPWR VPWR _12779_/D sky130_fd_sc_hd__clkbuf_1
X_06515_ _06515_/A _06527_/A VGND VGND VPWR VPWR _06520_/A sky130_fd_sc_hd__or2_1
XFILLER_22_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07495_ _08124_/A VGND VGND VPWR VPWR _07495_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09234_ _09234_/A VGND VGND VPWR VPWR _09234_/Y sky130_fd_sc_hd__inv_2
X_06446_ _06446_/A _06446_/B _06446_/C VGND VGND VPWR VPWR _06448_/B sky130_fd_sc_hd__and3_1
X_09165_ _09173_/A _09165_/B VGND VGND VPWR VPWR _09165_/Y sky130_fd_sc_hd__nand2_1
X_06377_ _13109_/D VGND VGND VPWR VPWR _06429_/A sky130_fd_sc_hd__inv_2
XFILLER_5_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08116_ _08161_/S _14005_/Q VGND VGND VPWR VPWR _08116_/X sky130_fd_sc_hd__or2b_1
XFILLER_147_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09096_ _09095_/B _09095_/C _09095_/A VGND VGND VPWR VPWR _09096_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_134_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08047_ _12961_/Q _13261_/Q _08051_/S VGND VGND VPWR VPWR _08048_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09998_ _10008_/S VGND VGND VPWR VPWR _10635_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08949_ _08978_/A _08978_/B VGND VGND VPWR VPWR _08951_/C sky130_fd_sc_hd__and2_1
XFILLER_29_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_68_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _13535_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11960_ _14297_/Q _11959_/X _11966_/S VGND VGND VPWR VPWR _11961_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10911_ _14745_/Q VGND VGND VPWR VPWR _11186_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11891_ _11891_/A VGND VGND VPWR VPWR _14242_/D sky130_fd_sc_hd__clkbuf_1
X_13630_ _14075_/CLK hold142/X VGND VGND VPWR VPWR _13630_/Q sky130_fd_sc_hd__dfxtp_1
X_10842_ _10842_/A VGND VGND VPWR VPWR _13181_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13561_ _13565_/CLK hold374/X VGND VGND VPWR VPWR _13561_/Q sky130_fd_sc_hd__dfxtp_1
X_10773_ _13008_/Q _10779_/B VGND VGND VPWR VPWR _10774_/A sky130_fd_sc_hd__and2_1
X_12512_ _12562_/S VGND VGND VPWR VPWR _12521_/S sky130_fd_sc_hd__buf_2
XFILLER_9_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13492_ _13722_/CLK hold218/X VGND VGND VPWR VPWR _13492_/Q sky130_fd_sc_hd__dfxtp_1
X_12443_ _12443_/A VGND VGND VPWR VPWR _14653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12374_ _12374_/A VGND VGND VPWR VPWR _14609_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14113_ _14605_/CLK hold26/X VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__dfxtp_1
X_11325_ _11325_/A VGND VGND VPWR VPWR _13768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14044_ _14050_/CLK _14044_/D VGND VGND VPWR VPWR _14044_/Q sky130_fd_sc_hd__dfxtp_1
X_11256_ _14036_/Q _14002_/Q _13842_/Q _14554_/Q _10993_/A _10995_/A VGND VGND VPWR
+ VPWR _11257_/A sky130_fd_sc_hd__mux4_1
XFILLER_125_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10207_ _10207_/A VGND VGND VPWR VPWR _14419_/D sky130_fd_sc_hd__clkbuf_1
X_11187_ _12584_/A VGND VGND VPWR VPWR _11187_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10138_ _10138_/A VGND VGND VPWR VPWR _14183_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_59_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _13076_/CLK sky130_fd_sc_hd__clkbuf_16
X_10069_ _14040_/D _10068_/X _14050_/D VGND VGND VPWR VPWR _10070_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13828_ _14709_/CLK _13828_/D VGND VGND VPWR VPWR _13828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13759_ _14707_/CLK _13759_/D VGND VGND VPWR VPWR _13759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06300_ _06300_/A VGND VGND VPWR VPWR _14184_/D sky130_fd_sc_hd__clkbuf_1
X_07280_ _07239_/X _07276_/X _07277_/Y _07279_/X VGND VGND VPWR VPWR _13133_/D sky130_fd_sc_hd__a31o_1
X_06231_ _06231_/A VGND VGND VPWR VPWR _06245_/B sky130_fd_sc_hd__clkbuf_1
X_06162_ _13855_/Q _06175_/B VGND VGND VPWR VPWR _06163_/A sky130_fd_sc_hd__and2_1
XFILLER_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold203 hold203/A VGND VGND VPWR VPWR hold203/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold214 hold214/A VGND VGND VPWR VPWR hold214/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold225 hold225/A VGND VGND VPWR VPWR hold225/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_06093_ _06093_/A VGND VGND VPWR VPWR _13937_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold236 hold236/A VGND VGND VPWR VPWR hold236/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_160_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold247 hold247/A VGND VGND VPWR VPWR hold247/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold258 hold258/A VGND VGND VPWR VPWR hold258/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold269 hold269/A VGND VGND VPWR VPWR hold269/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09921_ _09921_/A VGND VGND VPWR VPWR _12848_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ _13683_/Q _09851_/A _13684_/Q VGND VGND VPWR VPWR _09853_/C sky130_fd_sc_hd__a21o_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08803_ _13428_/Q VGND VGND VPWR VPWR _08851_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _09783_/A _09783_/B VGND VGND VPWR VPWR _09783_/Y sky130_fd_sc_hd__xnor2_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06995_ _13026_/Q _13027_/Q _06895_/B VGND VGND VPWR VPWR _07001_/B sky130_fd_sc_hd__o21ai_1
XFILLER_86_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08734_ _08724_/A _08728_/X _08741_/C _08733_/X VGND VGND VPWR VPWR _08734_/X sky130_fd_sc_hd__a31o_1
X_05946_ hold199/A _13862_/Q _13863_/Q _13866_/Q VGND VGND VPWR VPWR _05951_/C sky130_fd_sc_hd__and4_1
XFILLER_38_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08665_ _08665_/A _09472_/B VGND VGND VPWR VPWR _08665_/X sky130_fd_sc_hd__and2_1
XFILLER_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _13169_/D _07616_/B VGND VGND VPWR VPWR _07616_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _08596_/A _08596_/B VGND VGND VPWR VPWR _08605_/A sky130_fd_sc_hd__nor2_1
XFILLER_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07547_ _07547_/A _07547_/B VGND VGND VPWR VPWR _07548_/B sky130_fd_sc_hd__and2_1
XFILLER_22_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07478_ _13147_/Q _07579_/B _07477_/X VGND VGND VPWR VPWR _07488_/A sky130_fd_sc_hd__a21oi_1
XFILLER_139_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09217_ _13543_/Q _09228_/B VGND VGND VPWR VPWR _09226_/A sky130_fd_sc_hd__and2_1
X_06429_ _06429_/A _06429_/B _06429_/C VGND VGND VPWR VPWR _06429_/X sky130_fd_sc_hd__and3_1
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09148_ _09159_/A _09149_/B VGND VGND VPWR VPWR _09156_/B sky130_fd_sc_hd__or2_1
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09079_ _09079_/A VGND VGND VPWR VPWR _12772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11110_ _14307_/Q _14477_/Q _14233_/Q _14063_/Q _11066_/X _11067_/X VGND VGND VPWR
+ VPWR _11110_/X sky130_fd_sc_hd__mux4_1
X_12090_ _12090_/A VGND VGND VPWR VPWR _14462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11041_ _11041_/A _11013_/X VGND VGND VPWR VPWR _11041_/X sky130_fd_sc_hd__or2b_1
XFILLER_1_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12992_ _13351_/CLK _12992_/D VGND VGND VPWR VPWR hold154/A sky130_fd_sc_hd__dfxtp_2
XFILLER_18_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14731_ _14732_/CLK _14731_/D VGND VGND VPWR VPWR _14731_/Q sky130_fd_sc_hd__dfxtp_1
X_11943_ _11943_/A VGND VGND VPWR VPWR _14277_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _14717_/CLK _14662_/D VGND VGND VPWR VPWR _14662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ _11874_/A VGND VGND VPWR VPWR _14234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13613_ _13635_/CLK _13613_/D repeater57/X VGND VGND VPWR VPWR _13613_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10825_ _13132_/Q _10893_/A VGND VGND VPWR VPWR _10826_/A sky130_fd_sc_hd__and2_1
X_14593_ _14644_/CLK _14593_/D VGND VGND VPWR VPWR _14593_/Q sky130_fd_sc_hd__dfxtp_1
X_13544_ _13552_/CLK _13544_/D _12609_/A VGND VGND VPWR VPWR _13544_/Q sky130_fd_sc_hd__dfrtp_2
X_10756_ _10756_/A VGND VGND VPWR VPWR _13042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13475_ _13476_/CLK _13475_/D VGND VGND VPWR VPWR _13475_/Q sky130_fd_sc_hd__dfxtp_2
X_10687_ _12880_/Q _10687_/B VGND VGND VPWR VPWR _10688_/A sky130_fd_sc_hd__and2_1
X_12426_ _12484_/A _12484_/B input7/X VGND VGND VPWR VPWR _12427_/A sky130_fd_sc_hd__and3_1
XFILLER_127_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12357_ _12357_/A VGND VGND VPWR VPWR _14601_/D sky130_fd_sc_hd__clkbuf_1
X_11308_ _13763_/Q _11307_/X _11311_/S VGND VGND VPWR VPWR _11309_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12288_ _12288_/A VGND VGND VPWR VPWR _14560_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14027_ _14543_/CLK _14027_/D VGND VGND VPWR VPWR _14027_/Q sky130_fd_sc_hd__dfxtp_1
X_11239_ _14278_/Q _14669_/Q _13776_/Q _14724_/Q _10914_/A _10918_/A VGND VGND VPWR
+ VPWR _11240_/B sky130_fd_sc_hd__mux4_1
XFILLER_68_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06780_ _07861_/S VGND VGND VPWR VPWR _06793_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08450_ _08535_/A _08671_/B _08450_/C _08450_/D VGND VGND VPWR VPWR _08490_/A sky130_fd_sc_hd__nand4_2
XFILLER_17_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07401_ _07401_/A _07401_/B _07401_/C VGND VGND VPWR VPWR _07461_/C sky130_fd_sc_hd__or3_1
XFILLER_50_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08381_ _08381_/A VGND VGND VPWR VPWR _12723_/D sky130_fd_sc_hd__clkbuf_1
X_07332_ _13663_/Q _13661_/Q _13659_/Q _13657_/Q _07344_/S _07247_/X VGND VGND VPWR
+ VPWR _07333_/B sky130_fd_sc_hd__mux4_1
X_07263_ _07255_/B _07258_/B _07255_/A VGND VGND VPWR VPWR _07276_/A sky130_fd_sc_hd__o21ba_1
XFILLER_164_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14757__68 VGND VGND VPWR VPWR _14757__68/HI data_o[31] sky130_fd_sc_hd__conb_1
X_09002_ _09002_/A _09002_/B VGND VGND VPWR VPWR _09003_/B sky130_fd_sc_hd__xnor2_1
X_06214_ _14379_/Q _06215_/C _06215_/D _06216_/A VGND VGND VPWR VPWR _06324_/B sky130_fd_sc_hd__and4_1
XFILLER_164_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07194_ _07201_/A _07194_/B VGND VGND VPWR VPWR _07196_/C sky130_fd_sc_hd__xnor2_1
XFILLER_117_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06145_ _14162_/Q _06292_/A _06145_/C _06145_/D VGND VGND VPWR VPWR _06146_/B sky130_fd_sc_hd__or4_1
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06076_ _06076_/A _06076_/B VGND VGND VPWR VPWR _06076_/Y sky130_fd_sc_hd__nor2_1
XFILLER_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09904_ _09974_/S VGND VGND VPWR VPWR _09913_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_116_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09835_ _09835_/A VGND VGND VPWR VPWR _13681_/D sky130_fd_sc_hd__clkbuf_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09766_ _09778_/A _09778_/B _09768_/B VGND VGND VPWR VPWR _09769_/B sky130_fd_sc_hd__and3_1
X_06978_ _06978_/A _06978_/B VGND VGND VPWR VPWR _06979_/B sky130_fd_sc_hd__nand2_1
XFILLER_74_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08717_ _08689_/B _08715_/Y _08744_/A VGND VGND VPWR VPWR _08718_/B sky130_fd_sc_hd__a21oi_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05929_ _13716_/Q _13717_/Q _13718_/Q _13719_/Q VGND VGND VPWR VPWR _05935_/A sky130_fd_sc_hd__or4_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09697_ _09697_/A _09697_/B VGND VGND VPWR VPWR _09697_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_27_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _08650_/B VGND VGND VPWR VPWR _09464_/B sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08579_ _08635_/B _08444_/X _08579_/S VGND VGND VPWR VPWR _08579_/X sky130_fd_sc_hd__mux2_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10610_ _14040_/Q _14039_/Q _14042_/Q _14041_/Q VGND VGND VPWR VPWR _10610_/X sky130_fd_sc_hd__or4_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11590_ _11590_/A VGND VGND VPWR VPWR _13876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10541_ _10525_/A _10523_/Y _10533_/A _10509_/A VGND VGND VPWR VPWR _10542_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13260_ _13264_/CLK _13260_/D hold1/X VGND VGND VPWR VPWR _13260_/Q sky130_fd_sc_hd__dfrtp_1
X_10472_ _10463_/A _10463_/B _10466_/A VGND VGND VPWR VPWR _10480_/A sky130_fd_sc_hd__a21oi_1
XFILLER_136_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12211_ _12211_/A VGND VGND VPWR VPWR _14514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13191_ _13606_/CLK _13191_/D VGND VGND VPWR VPWR hold471/A sky130_fd_sc_hd__dfxtp_1
XFILLER_151_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12142_ _12142_/A VGND VGND VPWR VPWR _14485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12073_ _12073_/A VGND VGND VPWR VPWR _14454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11024_ _11166_/A VGND VGND VPWR VPWR _11024_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12975_ _13274_/CLK hold247/X VGND VGND VPWR VPWR _12975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14714_ _14714_/CLK _14714_/D VGND VGND VPWR VPWR _14714_/Q sky130_fd_sc_hd__dfxtp_1
X_11926_ _11926_/A VGND VGND VPWR VPWR _14269_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _14645_/CLK _14645_/D VGND VGND VPWR VPWR _14645_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _11857_/A VGND VGND VPWR VPWR _14226_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10808_ _13024_/Q _10812_/B VGND VGND VPWR VPWR _10809_/A sky130_fd_sc_hd__and2_1
X_14576_ _14615_/CLK _14576_/D VGND VGND VPWR VPWR _14576_/Q sky130_fd_sc_hd__dfxtp_1
X_11788_ _11788_/A VGND VGND VPWR VPWR _14087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13527_ _13528_/CLK _13527_/D _12609_/A VGND VGND VPWR VPWR _13527_/Q sky130_fd_sc_hd__dfrtp_1
X_10739_ _10739_/A VGND VGND VPWR VPWR _12946_/D sky130_fd_sc_hd__clkbuf_1
X_13458_ _13626_/CLK _13458_/D repeater57/X VGND VGND VPWR VPWR _13458_/Q sky130_fd_sc_hd__dfrtp_1
X_12409_ _12502_/B VGND VGND VPWR VPWR _12418_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_127_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13389_ _14690_/CLK _13389_/D VGND VGND VPWR VPWR _13389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07950_ _13268_/Q _13269_/Q _13270_/Q _13271_/Q _07989_/B VGND VGND VPWR VPWR _07975_/A
+ sky130_fd_sc_hd__o41a_1
X_06901_ _13015_/Q _07968_/B VGND VGND VPWR VPWR _06914_/A sky130_fd_sc_hd__nand2_1
X_07881_ _07881_/A _07881_/B _07892_/D VGND VGND VPWR VPWR _07881_/Y sky130_fd_sc_hd__nand3_1
XFILLER_96_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09620_ _13407_/Q _13605_/Q _09620_/S VGND VGND VPWR VPWR _09621_/A sky130_fd_sc_hd__mux2_1
X_06832_ _13010_/Q _07889_/B VGND VGND VPWR VPWR _06846_/A sky130_fd_sc_hd__nand2_1
XFILLER_96_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09551_ _09556_/A _09551_/B VGND VGND VPWR VPWR _09559_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06763_ _13032_/Q VGND VGND VPWR VPWR _07861_/S sky130_fd_sc_hd__clkbuf_2
X_08502_ _09388_/B _08500_/X _09404_/S VGND VGND VPWR VPWR _08503_/A sky130_fd_sc_hd__mux2_1
X_09482_ _13605_/Q _09530_/B VGND VGND VPWR VPWR _09484_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06694_ _06695_/B VGND VGND VPWR VPWR _07819_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08433_ _14255_/Q _14253_/Q _14251_/Q _14249_/Q _08472_/A _13475_/Q VGND VGND VPWR
+ VPWR _08564_/B sky130_fd_sc_hd__mux4_1
XFILLER_51_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08364_ _08397_/A VGND VGND VPWR VPWR _08373_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_149_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07315_ _13136_/Q _09112_/B VGND VGND VPWR VPWR _07316_/A sky130_fd_sc_hd__nand2_1
XFILLER_149_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08295_ _13370_/Q _08294_/A _13371_/Q VGND VGND VPWR VPWR _08296_/C sky130_fd_sc_hd__a21o_1
XFILLER_137_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07246_ _07344_/S _13390_/Q VGND VGND VPWR VPWR _07246_/X sky130_fd_sc_hd__and2b_1
XFILLER_152_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07177_ _07178_/A _07178_/B _07177_/C VGND VGND VPWR VPWR _07196_/A sky130_fd_sc_hd__or3_1
XFILLER_105_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06128_ _06126_/X _06122_/X _10106_/A VGND VGND VPWR VPWR _06129_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06059_ _06059_/A VGND VGND VPWR VPWR _13918_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09818_ _09818_/A VGND VGND VPWR VPWR _13679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09749_ _09749_/A _09749_/B VGND VGND VPWR VPWR _09753_/A sky130_fd_sc_hd__or2_2
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _13602_/CLK _12760_/D VGND VGND VPWR VPWR hold141/A sky130_fd_sc_hd__dfxtp_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _12662_/D _12661_/D _12662_/Q _11274_/Y VGND VGND VPWR VPWR _12564_/A sky130_fd_sc_hd__o31a_1
XFILLER_15_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _13303_/CLK _12691_/D VGND VGND VPWR VPWR hold418/A sky130_fd_sc_hd__dfxtp_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14430_ _14692_/CLK _14430_/D VGND VGND VPWR VPWR hold187/A sky130_fd_sc_hd__dfxtp_2
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _11642_/A VGND VGND VPWR VPWR _13996_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14361_ _14425_/CLK hold354/X VGND VGND VPWR VPWR _14361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11573_ _11573_/A VGND VGND VPWR VPWR _13868_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput18 data_i[30] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13312_ _14275_/CLK hold81/X VGND VGND VPWR VPWR _13312_/Q sky130_fd_sc_hd__dfxtp_1
Xinput29 rts_i VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__buf_4
X_10524_ _10512_/A _10509_/A _10533_/A _10523_/Y VGND VGND VPWR VPWR _10525_/B sky130_fd_sc_hd__a31o_1
XFILLER_128_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14292_ _14292_/CLK _14292_/D VGND VGND VPWR VPWR hold264/A sky130_fd_sc_hd__dfxtp_1
XFILLER_156_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13243_ _14702_/CLK _14702_/Q VGND VGND VPWR VPWR _13515_/D sky130_fd_sc_hd__dfxtp_2
X_10455_ _10441_/A _10485_/B _10456_/C VGND VGND VPWR VPWR _10461_/B sky130_fd_sc_hd__a21o_1
XFILLER_151_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13174_ _14012_/CLK _13174_/D VGND VGND VPWR VPWR hold360/A sky130_fd_sc_hd__dfxtp_1
X_10386_ _10386_/A _13518_/Q VGND VGND VPWR VPWR _10388_/A sky130_fd_sc_hd__nand2_1
X_12125_ _12125_/A VGND VGND VPWR VPWR _14477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12056_ _12056_/A VGND VGND VPWR VPWR _14446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11007_ _12566_/A VGND VGND VPWR VPWR _12645_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_38_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12958_ _13039_/CLK hold32/X VGND VGND VPWR VPWR _12958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11909_ _11931_/A VGND VGND VPWR VPWR _11918_/S sky130_fd_sc_hd__buf_2
XFILLER_34_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12889_ _12970_/CLK _12889_/D repeater59/X VGND VGND VPWR VPWR _12889_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14628_ _14690_/CLK _14628_/D VGND VGND VPWR VPWR _14628_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14559_ _14749_/CLK _14559_/D VGND VGND VPWR VPWR _14559_/Q sky130_fd_sc_hd__dfxtp_1
X_07100_ _07131_/A _07131_/B VGND VGND VPWR VPWR _07101_/B sky130_fd_sc_hd__xnor2_1
X_08080_ _12976_/Q _13276_/Q _08084_/S VGND VGND VPWR VPWR _08081_/A sky130_fd_sc_hd__mux2_1
X_07031_ _07031_/A _07141_/A VGND VGND VPWR VPWR _07032_/B sky130_fd_sc_hd__nand2_1
XFILLER_127_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08982_ _08989_/A _08982_/B VGND VGND VPWR VPWR _08984_/C sky130_fd_sc_hd__xnor2_1
XFILLER_103_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07933_ _06976_/X _07931_/X _07932_/X VGND VGND VPWR VPWR _13269_/D sky130_fd_sc_hd__a21o_1
XFILLER_130_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07864_ _06796_/A _07863_/C _13261_/Q VGND VGND VPWR VPWR _07885_/D sky130_fd_sc_hd__a21oi_1
XFILLER_68_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09603_ _13399_/Q _13597_/Q _09609_/S VGND VGND VPWR VPWR _09604_/A sky130_fd_sc_hd__mux2_2
X_06815_ _07863_/B _06813_/B _06813_/C _06800_/A VGND VGND VPWR VPWR _07878_/C sky130_fd_sc_hd__o22ai_4
X_07795_ _07745_/C _07788_/A _07785_/C _07785_/B VGND VGND VPWR VPWR _07796_/B sky130_fd_sc_hd__o211a_1
XFILLER_83_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09534_ _09534_/A _09534_/B _09534_/C _09532_/C VGND VGND VPWR VPWR _09535_/B sky130_fd_sc_hd__or4b_1
X_06746_ _13036_/Q _13353_/Q _06746_/S VGND VGND VPWR VPWR _06746_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09465_ _09475_/A _09465_/B VGND VGND VPWR VPWR _09477_/A sky130_fd_sc_hd__nand2_1
X_06677_ _06690_/A _06690_/B VGND VGND VPWR VPWR _07813_/B sky130_fd_sc_hd__xor2_1
XFILLER_51_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08416_ hold340/X _13384_/Q _08418_/S VGND VGND VPWR VPWR _08417_/A sky130_fd_sc_hd__mux2_1
X_09396_ _09396_/A _09419_/A _09419_/B VGND VGND VPWR VPWR _09396_/Y sky130_fd_sc_hd__nand3_1
XFILLER_138_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08347_ _10831_/A VGND VGND VPWR VPWR _10891_/B sky130_fd_sc_hd__buf_2
XFILLER_149_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08278_ _08278_/A VGND VGND VPWR VPWR _13368_/D sky130_fd_sc_hd__clkbuf_1
X_07229_ _13665_/Q _13663_/Q _13661_/Q _13659_/Q _13170_/Q _13171_/Q VGND VGND VPWR
+ VPWR _07361_/B sky130_fd_sc_hd__mux4_2
XFILLER_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10240_ _10240_/A VGND VGND VPWR VPWR _14529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10171_ _10171_/A VGND VGND VPWR VPWR _14135_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13930_ _13972_/CLK hold52/X VGND VGND VPWR VPWR hold498/A sky130_fd_sc_hd__dfxtp_1
XFILLER_75_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13861_ _14657_/CLK _13861_/D VGND VGND VPWR VPWR _13861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12812_ _13622_/CLK _12812_/D VGND VGND VPWR VPWR hold128/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13792_ _13799_/CLK _13792_/D VGND VGND VPWR VPWR _13792_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _14250_/CLK _12743_/D VGND VGND VPWR VPWR hold116/A sky130_fd_sc_hd__dfxtp_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _14647_/CLK _12674_/D VGND VGND VPWR VPWR hold119/A sky130_fd_sc_hd__dfxtp_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _14413_/CLK _14413_/D VGND VGND VPWR VPWR _14413_/Q sky130_fd_sc_hd__dfxtp_1
X_11625_ _11636_/A VGND VGND VPWR VPWR _11634_/S sky130_fd_sc_hd__buf_2
XFILLER_156_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14344_ _14357_/CLK hold106/X VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_155_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11556_ _11556_/A VGND VGND VPWR VPWR _13860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10507_ _14430_/D VGND VGND VPWR VPWR _10512_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14275_ _14275_/CLK _14275_/D VGND VGND VPWR VPWR _14275_/Q sky130_fd_sc_hd__dfxtp_1
X_11487_ _11487_/A VGND VGND VPWR VPWR _13830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13226_ _13605_/CLK hold246/X VGND VGND VPWR VPWR _13226_/Q sky130_fd_sc_hd__dfxtp_1
X_10438_ _10441_/A _10438_/B VGND VGND VPWR VPWR _14004_/D sky130_fd_sc_hd__nor2_1
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _13552_/CLK _13157_/D _12609_/A VGND VGND VPWR VPWR _13157_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10369_ _13518_/Q VGND VGND VPWR VPWR _10374_/A sky130_fd_sc_hd__clkbuf_2
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _12130_/A VGND VGND VPWR VPWR _12117_/S sky130_fd_sc_hd__clkbuf_2
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _13558_/CLK hold145/X VGND VGND VPWR VPWR _13088_/Q sky130_fd_sc_hd__dfxtp_1
X_12039_ _14367_/D _14369_/D _12039_/C _14382_/Q VGND VGND VPWR VPWR _12040_/A sky130_fd_sc_hd__or4b_1
XFILLER_78_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_1_0_clk clkbuf_4_1_0_clk/A VGND VGND VPWR VPWR clkbuf_4_1_0_clk/X sky130_fd_sc_hd__clkbuf_2
X_06600_ _12899_/Q _06597_/A _06599_/X VGND VGND VPWR VPWR _06601_/B sky130_fd_sc_hd__o21ai_1
X_07580_ _13161_/Q _09284_/B VGND VGND VPWR VPWR _07581_/B sky130_fd_sc_hd__nor2_1
XFILLER_92_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06531_ _06531_/A VGND VGND VPWR VPWR _12887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09250_ _13548_/Q _09250_/B VGND VGND VPWR VPWR _09255_/B sky130_fd_sc_hd__xor2_1
XFILLER_22_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06462_ _12881_/Q _06462_/B VGND VGND VPWR VPWR _06462_/X sky130_fd_sc_hd__or2_1
X_08201_ _13361_/Q _08201_/B VGND VGND VPWR VPWR _08202_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09181_ _09106_/X _09186_/B _09180_/Y _07445_/X VGND VGND VPWR VPWR _13537_/D sky130_fd_sc_hd__a31o_1
X_06393_ _12671_/Q _14438_/Q _14436_/Q _14434_/Q _06425_/S _13107_/D VGND VGND VPWR
+ VPWR _06504_/B sky130_fd_sc_hd__mux4_2
XFILLER_147_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08132_ _08164_/A _08152_/C VGND VGND VPWR VPWR _08135_/B sky130_fd_sc_hd__and2_1
XFILLER_147_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08063_ _08063_/A VGND VGND VPWR VPWR _12692_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07014_ hold425/A VGND VGND VPWR VPWR _07119_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08965_ _08966_/A _08966_/B _08965_/C VGND VGND VPWR VPWR _08984_/A sky130_fd_sc_hd__or3_1
XFILLER_75_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07916_ _07916_/A _07916_/B VGND VGND VPWR VPWR _07917_/B sky130_fd_sc_hd__nor2_1
XFILLER_29_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08896_ _13520_/D VGND VGND VPWR VPWR _08951_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07847_ _07847_/A _07859_/A VGND VGND VPWR VPWR _07858_/D sky130_fd_sc_hd__or2_2
XFILLER_29_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07778_ _07778_/A _07778_/B _07778_/C VGND VGND VPWR VPWR _07779_/B sky130_fd_sc_hd__and3_1
XFILLER_71_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09517_ _13610_/Q _09530_/B VGND VGND VPWR VPWR _09519_/A sky130_fd_sc_hd__nand2_1
X_06729_ _06729_/A VGND VGND VPWR VPWR _06730_/A sky130_fd_sc_hd__inv_2
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09448_ _09454_/B _09448_/B _09448_/C _09448_/D VGND VGND VPWR VPWR _09448_/Y sky130_fd_sc_hd__nor4_1
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09379_ _08784_/X _09377_/Y _09378_/X _08485_/X VGND VGND VPWR VPWR _13591_/D sky130_fd_sc_hd__a31o_1
XFILLER_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11410_ _13728_/Q _11416_/B VGND VGND VPWR VPWR _11411_/A sky130_fd_sc_hd__and2_1
X_12390_ _14617_/Q _12019_/X _12394_/S VGND VGND VPWR VPWR _12391_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11341_ _13888_/Q _13885_/Q _13889_/Q VGND VGND VPWR VPWR _11342_/C sky130_fd_sc_hd__a21o_1
XFILLER_4_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14060_ _14495_/CLK _14060_/D VGND VGND VPWR VPWR _14060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11272_ _14694_/Q VGND VGND VPWR VPWR _11272_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13011_ _13298_/CLK _13011_/D repeater59/X VGND VGND VPWR VPWR _13011_/Q sky130_fd_sc_hd__dfrtp_1
X_10223_ _10223_/A VGND VGND VPWR VPWR _14399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10154_ _14149_/Q _10143_/X _10150_/A VGND VGND VPWR VPWR _14284_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10085_ _10016_/A _10063_/X _10072_/X VGND VGND VPWR VPWR _10085_/X sky130_fd_sc_hd__a21o_1
XFILLER_59_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_47_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13913_ _14179_/CLK _13913_/D VGND VGND VPWR VPWR _13913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13844_ _14042_/CLK hold146/X VGND VGND VPWR VPWR _13844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13775_ _14724_/CLK _13775_/D VGND VGND VPWR VPWR _13775_/Q sky130_fd_sc_hd__dfxtp_1
X_10987_ _11035_/A _10987_/B VGND VGND VPWR VPWR _10987_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12726_ _13372_/CLK _12726_/D VGND VGND VPWR VPWR hold63/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12657_ _14555_/CLK hold198/X _12609_/A VGND VGND VPWR VPWR hold510/A sky130_fd_sc_hd__dfrtp_1
X_11608_ _13981_/Q _11456_/X _11612_/S VGND VGND VPWR VPWR _11609_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12588_ _12583_/X _12584_/Y _12585_/X _12586_/Y _12587_/X VGND VGND VPWR VPWR _12591_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_129_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14327_ _14327_/CLK hold140/X VGND VGND VPWR VPWR _14327_/Q sky130_fd_sc_hd__dfxtp_1
X_11539_ _13629_/Q _11541_/B VGND VGND VPWR VPWR _11540_/A sky130_fd_sc_hd__and2_1
Xhold407 hold407/A VGND VGND VPWR VPWR hold407/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold418 hold418/A VGND VGND VPWR VPWR hold418/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold429 hold429/A VGND VGND VPWR VPWR hold429/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_14258_ _14704_/CLK _14258_/D VGND VGND VPWR VPWR _14258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13209_ _13593_/CLK hold88/X VGND VGND VPWR VPWR _13209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ _14201_/CLK _14189_/D VGND VGND VPWR VPWR _14189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08748_/Y _08749_/X _08684_/X VGND VGND VPWR VPWR _13459_/D sky130_fd_sc_hd__a21o_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05962_ _13643_/Q _13644_/Q _13645_/Q _05962_/D VGND VGND VPWR VPWR _05963_/D sky130_fd_sc_hd__or4_1
X_07701_ _07701_/A _07701_/B _13114_/Q _13115_/Q VGND VGND VPWR VPWR _07732_/A sky130_fd_sc_hd__and4_1
XFILLER_39_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08681_ _09569_/B VGND VGND VPWR VPWR _08787_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_26_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07632_ _07610_/B _07614_/B _07610_/A VGND VGND VPWR VPWR _07633_/B sky130_fd_sc_hd__o21ba_1
XFILLER_26_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07563_ _07548_/A _07548_/B _07559_/Y _07562_/X VGND VGND VPWR VPWR _07578_/A sky130_fd_sc_hd__a31oi_2
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09302_ _13289_/Q _13527_/Q _09310_/S VGND VGND VPWR VPWR _09303_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06514_ _12886_/Q _06514_/B VGND VGND VPWR VPWR _06527_/A sky130_fd_sc_hd__nor2_1
XFILLER_34_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07494_ _07411_/X _07498_/B _07493_/Y _07486_/X VGND VGND VPWR VPWR _13149_/D sky130_fd_sc_hd__a31o_1
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09233_ _09226_/A _09226_/B _09229_/A _09228_/X _09241_/A VGND VGND VPWR VPWR _09234_/A
+ sky130_fd_sc_hd__o311a_1
X_06445_ _06442_/X _06443_/X _06444_/Y _06382_/X VGND VGND VPWR VPWR _06446_/C sky130_fd_sc_hd__o22a_1
X_09164_ _13535_/Q _09164_/B VGND VGND VPWR VPWR _09165_/B sky130_fd_sc_hd__or2_1
X_06376_ _10296_/B VGND VGND VPWR VPWR _14635_/D sky130_fd_sc_hd__inv_2
XFILLER_147_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08115_ _13424_/Q VGND VGND VPWR VPWR _08161_/S sky130_fd_sc_hd__clkbuf_2
X_09095_ _09095_/A _09095_/B _09095_/C VGND VGND VPWR VPWR _09095_/X sky130_fd_sc_hd__or3_1
X_08046_ _08046_/A VGND VGND VPWR VPWR _12684_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09997_ _14637_/Q _09997_/B VGND VGND VPWR VPWR _10008_/S sky130_fd_sc_hd__xnor2_1
XFILLER_131_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08948_ _08951_/B VGND VGND VPWR VPWR _08991_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08879_ _13515_/D _13432_/Q VGND VGND VPWR VPWR _08881_/C sky130_fd_sc_hd__nand2_1
XFILLER_91_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10910_ _11262_/A VGND VGND VPWR VPWR _12645_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11890_ _14242_/Q _11516_/X _11894_/S VGND VGND VPWR VPWR _11891_/A sky130_fd_sc_hd__mux2_1
X_10841_ _13139_/Q _10841_/B VGND VGND VPWR VPWR _10842_/A sky130_fd_sc_hd__and2_1
XFILLER_32_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13560_ _13562_/CLK hold178/X VGND VGND VPWR VPWR _13560_/Q sky130_fd_sc_hd__dfxtp_1
X_10772_ _10772_/A VGND VGND VPWR VPWR _13049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12511_ _12545_/A VGND VGND VPWR VPWR _12562_/S sky130_fd_sc_hd__buf_2
XFILLER_40_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13491_ _13722_/CLK hold169/X VGND VGND VPWR VPWR _13491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12442_ _14653_/Q _14699_/Q _12450_/S VGND VGND VPWR VPWR _12443_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12373_ _14609_/Q _11994_/X _12375_/S VGND VGND VPWR VPWR _12374_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14112_ _14693_/CLK hold38/X VGND VGND VPWR VPWR hold266/A sky130_fd_sc_hd__dfxtp_1
X_11324_ _13768_/Q _11323_/X _11327_/S VGND VGND VPWR VPWR _11325_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14043_ _14050_/CLK _14043_/D VGND VGND VPWR VPWR _14043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11255_ _14318_/Q _14488_/Q _14244_/Q _14074_/Q _11208_/X _11209_/X VGND VGND VPWR
+ VPWR _11255_/X sky130_fd_sc_hd__mux4_1
X_10206_ _06222_/X _06321_/X _10206_/S VGND VGND VPWR VPWR _10207_/A sky130_fd_sc_hd__mux2_1
X_11186_ _11186_/A VGND VGND VPWR VPWR _11186_/X sky130_fd_sc_hd__buf_2
XFILLER_122_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10137_ _13869_/Q _13853_/Q _10137_/S VGND VGND VPWR VPWR _10138_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10068_ _13921_/Q _10056_/X _10063_/A VGND VGND VPWR VPWR _10068_/X sky130_fd_sc_hd__a21o_1
XFILLER_85_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13827_ _14539_/CLK _13827_/D VGND VGND VPWR VPWR _13827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13758_ _14705_/CLK _13758_/D VGND VGND VPWR VPWR _13758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12709_ _14012_/CLK _12709_/D VGND VGND VPWR VPWR hold223/A sky130_fd_sc_hd__dfxtp_1
X_13689_ _13700_/CLK _13689_/D repeater57/X VGND VGND VPWR VPWR _13689_/Q sky130_fd_sc_hd__dfrtp_1
X_06230_ _06230_/A VGND VGND VPWR VPWR _14427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06161_ _06161_/A VGND VGND VPWR VPWR _06175_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold204 hold204/A VGND VGND VPWR VPWR hold204/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold215 hold215/A VGND VGND VPWR VPWR hold215/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06092_ _13791_/Q _06105_/B VGND VGND VPWR VPWR _06093_/A sky130_fd_sc_hd__and2_1
XFILLER_117_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold226 hold226/A VGND VGND VPWR VPWR hold226/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold237 hold237/A VGND VGND VPWR VPWR hold237/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold248 hold248/A VGND VGND VPWR VPWR hold248/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09920_ _13485_/Q _13674_/Q _09924_/S VGND VGND VPWR VPWR _09921_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold259 hold259/A VGND VGND VPWR VPWR hold259/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09851_ _09851_/A _09858_/D VGND VGND VPWR VPWR _09851_/X sky130_fd_sc_hd__and2_1
XFILLER_124_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08802_ _13516_/D VGND VGND VPWR VPWR _08907_/A sky130_fd_sc_hd__clkbuf_2
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09782_ _09781_/Y _09773_/B _09770_/A VGND VGND VPWR VPWR _09783_/B sky130_fd_sc_hd__a21oi_1
XFILLER_39_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06994_ _06945_/X _06992_/Y _06993_/X _06974_/X VGND VGND VPWR VPWR _13027_/D sky130_fd_sc_hd__a31o_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _08733_/A VGND VGND VPWR VPWR _08733_/X sky130_fd_sc_hd__clkbuf_2
X_05945_ _13864_/Q _13865_/Q _05945_/C _05945_/D VGND VGND VPWR VPWR _05952_/A sky130_fd_sc_hd__nor4_1
XFILLER_67_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08664_ _08664_/A _08664_/B _08664_/C VGND VGND VPWR VPWR _08664_/Y sky130_fd_sc_hd__nand3_1
XFILLER_38_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07615_ _07620_/A _07620_/B VGND VGND VPWR VPWR _07616_/B sky130_fd_sc_hd__xnor2_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _08657_/A _08595_/B VGND VGND VPWR VPWR _08596_/B sky130_fd_sc_hd__nor2_1
XFILLER_41_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07546_ _13155_/Q _13156_/Q _09284_/B VGND VGND VPWR VPWR _07553_/B sky130_fd_sc_hd__o21ai_1
XFILLER_22_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07477_ _07504_/A _07477_/B VGND VGND VPWR VPWR _07477_/X sky130_fd_sc_hd__and2b_1
X_09216_ _09182_/X _09213_/X _09214_/Y _09215_/X VGND VGND VPWR VPWR _13542_/D sky130_fd_sc_hd__a31o_1
X_06428_ _14434_/Q _14432_/Q _06458_/S VGND VGND VPWR VPWR _06429_/C sky130_fd_sc_hd__mux2_1
XFILLER_5_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09147_ _09137_/Y _09146_/X _09161_/C VGND VGND VPWR VPWR _09149_/B sky130_fd_sc_hd__o21bai_1
XFILLER_136_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06359_ _06357_/Y _06358_/X _12875_/D VGND VGND VPWR VPWR _06360_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09078_ _13236_/Q _13465_/Q _09587_/S VGND VGND VPWR VPWR _09079_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08029_ _08029_/A VGND VGND VPWR VPWR _12674_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11040_ _14020_/Q _13986_/Q _13826_/Q _14538_/Q _11010_/X _11011_/X VGND VGND VPWR
+ VPWR _11041_/A sky130_fd_sc_hd__mux4_1
XFILLER_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12991_ _13351_/CLK _12991_/D VGND VGND VPWR VPWR hold177/A sky130_fd_sc_hd__dfxtp_1
X_11942_ _14277_/Q _11513_/X _11948_/S VGND VGND VPWR VPWR _11943_/A sky130_fd_sc_hd__mux2_1
X_14730_ _14732_/CLK _14730_/D VGND VGND VPWR VPWR _14730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _14716_/CLK _14661_/D VGND VGND VPWR VPWR _14661_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _14234_/Q _11491_/X _11875_/S VGND VGND VPWR VPWR _11874_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13612_ _13619_/CLK _13612_/D repeater57/X VGND VGND VPWR VPWR _13612_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ _10824_/A VGND VGND VPWR VPWR _13173_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _14644_/CLK _14592_/D VGND VGND VPWR VPWR _14592_/Q sky130_fd_sc_hd__dfxtp_1
X_13543_ _13562_/CLK _13543_/D _12609_/A VGND VGND VPWR VPWR _13543_/Q sky130_fd_sc_hd__dfrtp_2
X_10755_ _13000_/Q _10820_/A VGND VGND VPWR VPWR _10756_/A sky130_fd_sc_hd__and2_1
XFILLER_13_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13474_ _13476_/CLK _13474_/D VGND VGND VPWR VPWR _13474_/Q sky130_fd_sc_hd__dfxtp_1
X_10686_ _10686_/A VGND VGND VPWR VPWR _12922_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12425_ _12425_/A VGND VGND VPWR VPWR _14645_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_12356_ _14601_/Q _11968_/X _12364_/S VGND VGND VPWR VPWR _12357_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11307_ _14513_/Q VGND VGND VPWR VPWR _11307_/X sky130_fd_sc_hd__buf_2
X_12287_ _14560_/Q _11959_/X _12291_/S VGND VGND VPWR VPWR _12288_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14026_ _14713_/CLK _14026_/D VGND VGND VPWR VPWR _14026_/Q sky130_fd_sc_hd__dfxtp_1
X_11238_ _11238_/A VGND VGND VPWR VPWR _11238_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11169_ _13333_/Q _11150_/X _11158_/X _11168_/Y VGND VGND VPWR VPWR _13333_/D sky130_fd_sc_hd__o22a_1
XFILLER_68_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07400_ _07400_/A _07400_/B VGND VGND VPWR VPWR _07401_/C sky130_fd_sc_hd__nor2_2
XFILLER_90_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08380_ _13087_/Q _13368_/Q _08384_/S VGND VGND VPWR VPWR _08381_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07331_ _13172_/Q VGND VGND VPWR VPWR _07387_/A sky130_fd_sc_hd__inv_2
XFILLER_149_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07262_ _07239_/X _07257_/X _07258_/Y _07261_/X VGND VGND VPWR VPWR _13132_/D sky130_fd_sc_hd__a31o_1
XFILLER_137_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09001_ _08951_/C _08994_/A _08991_/C _08991_/B VGND VGND VPWR VPWR _09002_/B sky130_fd_sc_hd__o211a_1
X_06213_ _14407_/Q _14399_/Q _06321_/S VGND VGND VPWR VPWR _06216_/A sky130_fd_sc_hd__mux2_1
X_07193_ _07205_/A _07205_/B _07178_/A VGND VGND VPWR VPWR _07194_/B sky130_fd_sc_hd__a21oi_1
XFILLER_118_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06144_ _14162_/Q _06145_/C _06145_/D _06146_/A VGND VGND VPWR VPWR _06292_/B sky130_fd_sc_hd__and4_1
XFILLER_145_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06075_ hold498/A _06259_/A _06075_/C _06075_/D VGND VGND VPWR VPWR _06076_/B sky130_fd_sc_hd__or4_1
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09903_ _13700_/Q VGND VGND VPWR VPWR _09974_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_104_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09834_ _09829_/B _09833_/Y _09834_/S VGND VGND VPWR VPWR _09835_/A sky130_fd_sc_hd__mux2_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _09765_/A VGND VGND VPWR VPWR _13674_/D sky130_fd_sc_hd__clkbuf_1
X_06977_ _13025_/Q _08001_/B VGND VGND VPWR VPWR _06981_/B sky130_fd_sc_hd__xnor2_1
XFILLER_27_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08716_ _13451_/Q _13452_/Q _13453_/Q _13454_/Q _09550_/B VGND VGND VPWR VPWR _08744_/A
+ sky130_fd_sc_hd__o41a_1
X_05928_ _05928_/A _05928_/B _05928_/C VGND VGND VPWR VPWR _05928_/X sky130_fd_sc_hd__and3_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09696_ _09696_/A _09696_/B VGND VGND VPWR VPWR _09697_/B sky130_fd_sc_hd__nand2_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08647_ _08591_/A _08596_/B _08607_/C _08646_/Y _08566_/B VGND VGND VPWR VPWR _08650_/B
+ sky130_fd_sc_hd__o311a_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08578_ _08578_/A VGND VGND VPWR VPWR _08657_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07529_ _07530_/A _07530_/B _07530_/C VGND VGND VPWR VPWR _07529_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_23_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10540_ _10540_/A _10539_/X VGND VGND VPWR VPWR _10542_/A sky130_fd_sc_hd__or2b_1
XFILLER_22_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10471_ _10471_/A _10471_/B VGND VGND VPWR VPWR _14008_/D sky130_fd_sc_hd__xnor2_1
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12210_ _12215_/C _12222_/B _12210_/C VGND VGND VPWR VPWR _12211_/A sky130_fd_sc_hd__and3b_1
XFILLER_109_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13190_ _13423_/CLK _13190_/D VGND VGND VPWR VPWR hold147/A sky130_fd_sc_hd__dfxtp_1
XFILLER_124_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12141_ _14485_/Q _12016_/X _12147_/S VGND VGND VPWR VPWR _12142_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12072_ _11323_/X _14454_/Q _12074_/S VGND VGND VPWR VPWR _12073_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11023_ _11035_/A _11023_/B VGND VGND VPWR VPWR _11023_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12974_ _12974_/CLK hold302/X VGND VGND VPWR VPWR _12974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14713_ _14713_/CLK _14713_/D VGND VGND VPWR VPWR _14713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11925_ _14269_/Q _11488_/X _11929_/S VGND VGND VPWR VPWR _11926_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14644_ _14644_/CLK _14644_/D VGND VGND VPWR VPWR _14644_/Q sky130_fd_sc_hd__dfxtp_1
X_11856_ _14226_/Q _11465_/X _11864_/S VGND VGND VPWR VPWR _11857_/A sky130_fd_sc_hd__mux2_1
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10807_ _10807_/A VGND VGND VPWR VPWR _13065_/D sky130_fd_sc_hd__clkbuf_1
X_14575_ _14615_/CLK _14575_/D VGND VGND VPWR VPWR _14575_/Q sky130_fd_sc_hd__dfxtp_1
X_11787_ _13565_/Q _11795_/B VGND VGND VPWR VPWR _11788_/A sky130_fd_sc_hd__and2_1
XFILLER_158_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10738_ _12903_/Q _10742_/B VGND VGND VPWR VPWR _10739_/A sky130_fd_sc_hd__and2_1
X_13526_ _13528_/CLK _13526_/D _12609_/A VGND VGND VPWR VPWR _13526_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_159_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13457_ _13605_/CLK _13457_/D repeater57/X VGND VGND VPWR VPWR _13457_/Q sky130_fd_sc_hd__dfrtp_1
X_10669_ _14341_/Q _10671_/C _10656_/X VGND VGND VPWR VPWR _10669_/Y sky130_fd_sc_hd__o21ai_1
X_12408_ input29/X VGND VGND VPWR VPWR _12502_/B sky130_fd_sc_hd__buf_2
X_13388_ _14647_/CLK _13388_/D VGND VGND VPWR VPWR _13388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12339_ _12339_/A VGND VGND VPWR VPWR _14593_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06900_ _06899_/Y _06924_/A _06887_/A VGND VGND VPWR VPWR _06909_/A sky130_fd_sc_hd__o21a_1
XFILLER_96_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14009_ _14012_/CLK _14009_/D VGND VGND VPWR VPWR _14009_/Q sky130_fd_sc_hd__dfxtp_1
X_07880_ _07881_/A _07881_/B _07892_/D VGND VGND VPWR VPWR _07880_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06831_ _06863_/A _06829_/X _06840_/A VGND VGND VPWR VPWR _07889_/B sky130_fd_sc_hd__o21a_2
XFILLER_56_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09550_ _13615_/Q _09550_/B VGND VGND VPWR VPWR _09551_/B sky130_fd_sc_hd__or2_1
X_06762_ _06762_/A _06762_/B VGND VGND VPWR VPWR _06762_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_37_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08501_ _09422_/S VGND VGND VPWR VPWR _09404_/S sky130_fd_sc_hd__buf_2
X_09481_ _09475_/A _09473_/B _09478_/Y _09460_/B _09480_/Y VGND VGND VPWR VPWR _09510_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_64_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06693_ _06719_/A _06696_/B VGND VGND VPWR VPWR _06695_/B sky130_fd_sc_hd__and2b_1
XFILLER_51_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08432_ _13474_/Q VGND VGND VPWR VPWR _08472_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08363_ _08363_/A VGND VGND VPWR VPWR _12715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07314_ _09112_/B VGND VGND VPWR VPWR _09120_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_08294_ _08294_/A _08301_/D VGND VGND VPWR VPWR _08294_/X sky130_fd_sc_hd__and2_1
XFILLER_109_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07245_ _13170_/Q VGND VGND VPWR VPWR _07344_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_118_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07176_ _07150_/A _07150_/B _07175_/X VGND VGND VPWR VPWR _07177_/C sky130_fd_sc_hd__a21oi_1
XFILLER_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06127_ _06127_/A VGND VGND VPWR VPWR _10106_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_132_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06058_ _06056_/X _06052_/X _10019_/A VGND VGND VPWR VPWR _06059_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09817_ _09811_/B _09816_/Y _09834_/S VGND VGND VPWR VPWR _09818_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09748_ _13673_/Q _09748_/B VGND VGND VPWR VPWR _09749_/B sky130_fd_sc_hd__nor2_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _09720_/A _13668_/Q _09679_/C VGND VGND VPWR VPWR _09681_/A sky130_fd_sc_hd__and3_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11841_/A VGND VGND VPWR VPWR _12619_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _13303_/CLK _12690_/D VGND VGND VPWR VPWR hold459/A sky130_fd_sc_hd__dfxtp_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11641_ _13996_/Q _11504_/X _11645_/S VGND VGND VPWR VPWR _11642_/A sky130_fd_sc_hd__mux2_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14360_ _14536_/CLK _14360_/D VGND VGND VPWR VPWR _14360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11572_ _13644_/Q _11574_/B VGND VGND VPWR VPWR _11573_/A sky130_fd_sc_hd__and2_1
XFILLER_11_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13311_ _14275_/CLK hold448/X VGND VGND VPWR VPWR _13311_/Q sky130_fd_sc_hd__dfxtp_1
Xinput19 data_i[31] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__buf_2
XFILLER_156_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10523_ _10509_/A _10519_/A _10557_/A VGND VGND VPWR VPWR _10523_/Y sky130_fd_sc_hd__o21ai_1
X_14291_ _14292_/CLK hold283/X VGND VGND VPWR VPWR _14291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13242_ _14010_/CLK _13242_/D VGND VGND VPWR VPWR _13514_/D sky130_fd_sc_hd__dfxtp_1
X_10454_ hold62/A VGND VGND VPWR VPWR _10485_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13173_ _14012_/CLK _13173_/D VGND VGND VPWR VPWR hold224/A sky130_fd_sc_hd__dfxtp_1
XFILLER_163_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10385_ _13518_/Q _10382_/X _10405_/A VGND VGND VPWR VPWR _10390_/A sky130_fd_sc_hd__o21ba_1
XFILLER_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12124_ _14477_/Q _11991_/X _12128_/S VGND VGND VPWR VPWR _12125_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12055_ _11297_/X _14446_/Q _12063_/S VGND VGND VPWR VPWR _12056_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11006_ _13322_/Q _10907_/X _10999_/X _11005_/Y VGND VGND VPWR VPWR _13322_/D sky130_fd_sc_hd__o22a_1
XFILLER_19_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12957_ _13263_/CLK hold275/X VGND VGND VPWR VPWR _12957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11908_ _11908_/A VGND VGND VPWR VPWR _14261_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _12930_/CLK _12888_/D hold1/X VGND VGND VPWR VPWR _12888_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14627_ _14647_/CLK hold461/X VGND VGND VPWR VPWR _14627_/Q sky130_fd_sc_hd__dfxtp_1
X_11839_ _14150_/D _14152_/D _11839_/C _14165_/Q VGND VGND VPWR VPWR _11840_/A sky130_fd_sc_hd__or4b_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14558_ _14749_/CLK _14558_/D VGND VGND VPWR VPWR _14558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13509_ _13698_/CLK hold33/X VGND VGND VPWR VPWR _13509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14489_ _14749_/CLK _14489_/D VGND VGND VPWR VPWR _14489_/Q sky130_fd_sc_hd__dfxtp_1
X_07030_ _07086_/C VGND VGND VPWR VPWR _07141_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08981_ _08993_/A _08993_/B _08966_/A VGND VGND VPWR VPWR _08982_/B sky130_fd_sc_hd__a21oi_1
XFILLER_130_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07932_ _07932_/A VGND VGND VPWR VPWR _07932_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07863_ _13261_/Q _07863_/B _07863_/C VGND VGND VPWR VPWR _07885_/C sky130_fd_sc_hd__and3_1
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09602_ _09602_/A VGND VGND VPWR VPWR _12815_/D sky130_fd_sc_hd__clkbuf_1
X_06814_ _06881_/C VGND VGND VPWR VPWR _07878_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_07794_ _07789_/A _07788_/B _07790_/B _07790_/A VGND VGND VPWR VPWR _07797_/A sky130_fd_sc_hd__a22o_1
X_09533_ _09502_/X _09531_/Y _09532_/X _09506_/X VGND VGND VPWR VPWR _13612_/D sky130_fd_sc_hd__a31o_1
X_06745_ _06745_/A VGND VGND VPWR VPWR _06745_/X sky130_fd_sc_hd__clkbuf_2
X_09464_ _13603_/Q _09464_/B VGND VGND VPWR VPWR _09465_/B sky130_fd_sc_hd__or2_1
X_06676_ _06636_/Y _06799_/B _06675_/X _06634_/X VGND VGND VPWR VPWR _06690_/B sky130_fd_sc_hd__a22oi_4
XFILLER_12_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08415_ _08415_/A VGND VGND VPWR VPWR _12738_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09395_ _13594_/Q _09401_/B VGND VGND VPWR VPWR _09419_/B sky130_fd_sc_hd__xnor2_1
XFILLER_51_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08346_ _13468_/D VGND VGND VPWR VPWR _10831_/A sky130_fd_sc_hd__buf_4
XFILLER_20_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08277_ _08272_/B _08276_/Y _08286_/S VGND VGND VPWR VPWR _08278_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07228_ _13167_/Q _13172_/Q VGND VGND VPWR VPWR _07228_/X sky130_fd_sc_hd__and2b_1
XFILLER_152_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07159_ _07151_/A _07151_/B _07152_/A VGND VGND VPWR VPWR _07182_/A sky130_fd_sc_hd__a21o_1
XFILLER_152_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10170_ _10165_/X _10169_/X _14292_/D VGND VGND VPWR VPWR _10171_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13860_ _14656_/CLK _13860_/D VGND VGND VPWR VPWR _13860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12811_ _13635_/CLK _12811_/D VGND VGND VPWR VPWR hold385/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13791_ _13843_/CLK _13791_/D VGND VGND VPWR VPWR _13791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _14250_/CLK _12742_/D VGND VGND VPWR VPWR hold209/A sky130_fd_sc_hd__dfxtp_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _13525_/CLK _12673_/D VGND VGND VPWR VPWR hold257/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_190_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _14724_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11624_ _11624_/A VGND VGND VPWR VPWR _13988_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _14413_/CLK _14412_/D VGND VGND VPWR VPWR _14412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14343_ _14697_/CLK hold474/X VGND VGND VPWR VPWR _14343_/Q sky130_fd_sc_hd__dfxtp_1
X_11555_ _13636_/Q _11563_/B VGND VGND VPWR VPWR _11556_/A sky130_fd_sc_hd__and2_1
XFILLER_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10506_ _12990_/D VGND VGND VPWR VPWR _10521_/B sky130_fd_sc_hd__inv_2
XFILLER_156_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14274_ _14275_/CLK _14274_/D VGND VGND VPWR VPWR _14274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11486_ _13830_/Q _11485_/X _11495_/S VGND VGND VPWR VPWR _11487_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13225_ _13605_/CLK hold509/X VGND VGND VPWR VPWR _13225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10437_ hold186/A VGND VGND VPWR VPWR _10438_/B sky130_fd_sc_hd__inv_2
XFILLER_152_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13156_ _14530_/CLK _13156_/D _12609_/A VGND VGND VPWR VPWR _13156_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10368_ _13516_/Q VGND VGND VPWR VPWR _10432_/B sky130_fd_sc_hd__inv_2
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _12107_/A VGND VGND VPWR VPWR _14469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _13423_/CLK hold124/X VGND VGND VPWR VPWR _13087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10299_ _10299_/A VGND VGND VPWR VPWR _14585_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12038_ _14365_/D _14366_/D _14368_/D _14370_/D VGND VGND VPWR VPWR _12039_/C sky130_fd_sc_hd__or4_1
XFILLER_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13989_ _14713_/CLK _13989_/D VGND VGND VPWR VPWR _13989_/Q sky130_fd_sc_hd__dfxtp_1
X_06530_ _06525_/B _06529_/Y _06530_/S VGND VGND VPWR VPWR _06531_/A sky130_fd_sc_hd__mux2_1
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06461_ _12881_/Q _06462_/B VGND VGND VPWR VPWR _06463_/A sky130_fd_sc_hd__and2_1
XFILLER_22_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_181_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _14533_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08200_ _13361_/Q _08201_/B VGND VGND VPWR VPWR _08202_/A sky130_fd_sc_hd__and2_1
X_09180_ _09189_/A _09180_/B VGND VGND VPWR VPWR _09180_/Y sky130_fd_sc_hd__nand2_1
X_06392_ _06392_/A VGND VGND VPWR VPWR _10346_/A sky130_fd_sc_hd__clkbuf_2
X_08131_ _08126_/X _08270_/B _08128_/X _08129_/X _08228_/S _08162_/B VGND VGND VPWR
+ VPWR _08152_/C sky130_fd_sc_hd__mux4_1
XFILLER_30_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08062_ _12968_/Q _13268_/Q _08062_/S VGND VGND VPWR VPWR _08063_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07013_ _13036_/D _07013_/B VGND VGND VPWR VPWR _10647_/B sky130_fd_sc_hd__xnor2_1
XFILLER_134_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08964_ _08938_/A _08938_/B _08963_/X VGND VGND VPWR VPWR _08965_/C sky130_fd_sc_hd__a21oi_1
XFILLER_97_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07915_ _07909_/X _07913_/X _07914_/Y _06871_/X VGND VGND VPWR VPWR _13267_/D sky130_fd_sc_hd__a31o_1
X_08895_ _08895_/A _08895_/B _08895_/C VGND VGND VPWR VPWR _08911_/B sky130_fd_sc_hd__or3_1
XFILLER_68_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07846_ _13259_/Q _07846_/B _07846_/C VGND VGND VPWR VPWR _07859_/A sky130_fd_sc_hd__and3_1
XFILLER_57_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07777_ _07778_/A _07778_/B _07778_/C VGND VGND VPWR VPWR _07779_/A sky130_fd_sc_hd__a21oi_1
XFILLER_37_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09516_ _09514_/X _09515_/Y _09493_/X VGND VGND VPWR VPWR _13609_/D sky130_fd_sc_hd__a21o_1
X_06728_ _13002_/Q _07832_/B VGND VGND VPWR VPWR _06729_/A sky130_fd_sc_hd__and2_1
XFILLER_140_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09447_ _09447_/A _09447_/B _09447_/C _09447_/D VGND VGND VPWR VPWR _09448_/B sky130_fd_sc_hd__or4_1
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06659_ _06659_/A _06659_/B VGND VGND VPWR VPWR _06661_/A sky130_fd_sc_hd__or2_1
XFILLER_25_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_172_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _14492_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09378_ _09377_/B _09377_/C _09377_/A VGND VGND VPWR VPWR _09378_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08329_ _08329_/A VGND VGND VPWR VPWR _13380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11340_ _13888_/Q _13885_/Q _13889_/Q VGND VGND VPWR VPWR _11351_/C sky130_fd_sc_hd__and3_1
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11271_ _11271_/A VGND VGND VPWR VPWR _13750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13010_ _13298_/CLK _13010_/D repeater59/X VGND VGND VPWR VPWR _13010_/Q sky130_fd_sc_hd__dfrtp_1
X_10222_ _14100_/Q _14084_/Q _10224_/S VGND VGND VPWR VPWR _10223_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10153_ _10153_/A VGND VGND VPWR VPWR _14290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10084_ _10084_/A VGND VGND VPWR VPWR _13903_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_13912_ _14179_/CLK _13965_/Q VGND VGND VPWR VPWR _13912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13843_ _13843_/CLK _13843_/D VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__dfxtp_2
XFILLER_90_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10986_ _14260_/Q _14651_/Q _13758_/Q _14706_/Q _10940_/X _10942_/X VGND VGND VPWR
+ VPWR _10987_/B sky130_fd_sc_hd__mux4_1
X_13774_ _14722_/CLK _13774_/D VGND VGND VPWR VPWR _13774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12725_ _13606_/CLK _12725_/D VGND VGND VPWR VPWR hold444/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_163_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _14530_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_130_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12656_ _14082_/CLK hold512/X _12609_/A VGND VGND VPWR VPWR hold198/A sky130_fd_sc_hd__dfrtp_1
XFILLER_90_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11607_ _11607_/A VGND VGND VPWR VPWR _13980_/D sky130_fd_sc_hd__clkbuf_1
X_12587_ _14748_/Q _14733_/Q VGND VGND VPWR VPWR _12587_/X sky130_fd_sc_hd__xor2_1
XFILLER_157_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14326_ _14688_/CLK _14326_/D VGND VGND VPWR VPWR _14326_/Q sky130_fd_sc_hd__dfxtp_1
X_11538_ _11538_/A VGND VGND VPWR VPWR _13852_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold408 hold408/A VGND VGND VPWR VPWR hold408/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold419 hold419/A VGND VGND VPWR VPWR hold419/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_11469_ _14700_/Q VGND VGND VPWR VPWR _11469_/X sky130_fd_sc_hd__clkbuf_2
X_14257_ _14533_/CLK _14257_/D VGND VGND VPWR VPWR _14257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13208_ _13593_/CLK hold65/X VGND VGND VPWR VPWR _13208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14188_ _14201_/CLK _14188_/D VGND VGND VPWR VPWR _14188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13139_ _13434_/CLK _13139_/D repeater56/X VGND VGND VPWR VPWR _13139_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05961_ _13635_/Q _13636_/Q _13637_/Q _13642_/Q VGND VGND VPWR VPWR _05962_/D sky130_fd_sc_hd__or4_1
XFILLER_97_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07700_ _07721_/A _07772_/B _07772_/D _07701_/A VGND VGND VPWR VPWR _07702_/A sky130_fd_sc_hd__a22oi_1
XFILLER_94_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08680_ _09562_/B VGND VGND VPWR VPWR _09569_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_07631_ _07641_/A _07631_/B VGND VGND VPWR VPWR _07640_/B sky130_fd_sc_hd__xnor2_1
XFILLER_66_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07562_ _13155_/Q _13156_/Q _13157_/Q _13158_/Q _09271_/B VGND VGND VPWR VPWR _07562_/X
+ sky130_fd_sc_hd__o41a_1
X_09301_ _09323_/A VGND VGND VPWR VPWR _09310_/S sky130_fd_sc_hd__clkbuf_2
X_06513_ _12886_/Q _06513_/B _06563_/B VGND VGND VPWR VPWR _06515_/A sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_154_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _14709_/CLK sky130_fd_sc_hd__clkbuf_16
X_07493_ _07493_/A _07493_/B _07504_/C VGND VGND VPWR VPWR _07493_/Y sky130_fd_sc_hd__nand3_1
X_09232_ _13545_/Q _09237_/B VGND VGND VPWR VPWR _09241_/A sky130_fd_sc_hd__xor2_1
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06444_ _06444_/A _06455_/A VGND VGND VPWR VPWR _06444_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09163_ _13535_/Q _09163_/B VGND VGND VPWR VPWR _09173_/A sky130_fd_sc_hd__nand2_1
X_06375_ hold118/X _10293_/A VGND VGND VPWR VPWR _10296_/B sky130_fd_sc_hd__nand2_1
X_08114_ _08143_/A _13426_/Q VGND VGND VPWR VPWR _08114_/X sky130_fd_sc_hd__or2b_1
X_09094_ _13525_/Q _09101_/B VGND VGND VPWR VPWR _09095_/C sky130_fd_sc_hd__and2_1
XFILLER_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08045_ _12960_/Q _13260_/Q _08051_/S VGND VGND VPWR VPWR _08046_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09996_ _13389_/Q _14628_/Q _14647_/Q VGND VGND VPWR VPWR _09997_/B sky130_fd_sc_hd__mux2_1
XFILLER_131_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08947_ _08939_/A _08939_/B _08940_/A VGND VGND VPWR VPWR _08970_/A sky130_fd_sc_hd__a21o_1
X_08878_ _13516_/D _13517_/D _08929_/B _13431_/Q VGND VGND VPWR VPWR _08881_/B sky130_fd_sc_hd__and4_2
XFILLER_151_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07829_ _07833_/B _07829_/B VGND VGND VPWR VPWR _07829_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_38_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10840_ _10840_/A VGND VGND VPWR VPWR _13180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10771_ _13007_/Q _10779_/B VGND VGND VPWR VPWR _10772_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_145_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _14610_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12510_ _12510_/A _12041_/C VGND VGND VPWR VPWR _12545_/A sky130_fd_sc_hd__or2b_4
X_13490_ _13722_/CLK hold129/X VGND VGND VPWR VPWR _13490_/Q sky130_fd_sc_hd__dfxtp_1
X_12441_ _12463_/A VGND VGND VPWR VPWR _12450_/S sky130_fd_sc_hd__buf_2
XFILLER_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12372_ _12372_/A VGND VGND VPWR VPWR _14608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14111_ _14693_/CLK hold266/X VGND VGND VPWR VPWR hold87/A sky130_fd_sc_hd__dfxtp_1
X_11323_ _14518_/Q VGND VGND VPWR VPWR _11323_/X sky130_fd_sc_hd__buf_2
Xclkbuf_4_0_0_clk clkbuf_4_1_0_clk/A VGND VGND VPWR VPWR clkbuf_4_0_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11254_ _13340_/Q _10962_/A _11247_/X _11253_/Y VGND VGND VPWR VPWR _13340_/D sky130_fd_sc_hd__o22a_1
X_14042_ _14042_/CLK _14042_/D VGND VGND VPWR VPWR _14042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10205_ _10205_/A VGND VGND VPWR VPWR _14418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11185_ _11185_/A VGND VGND VPWR VPWR _11242_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10136_ _10136_/A VGND VGND VPWR VPWR _14182_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10067_ _13917_/Q _10056_/X _10063_/A VGND VGND VPWR VPWR _14040_/D sky130_fd_sc_hd__a21o_1
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13826_ _14697_/CLK _13826_/D VGND VGND VPWR VPWR _13826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_136_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _14047_/CLK sky130_fd_sc_hd__clkbuf_16
X_13757_ _14705_/CLK _13757_/D VGND VGND VPWR VPWR _13757_/Q sky130_fd_sc_hd__dfxtp_1
X_10969_ _11186_/A VGND VGND VPWR VPWR _10969_/X sky130_fd_sc_hd__clkbuf_4
X_12708_ _13565_/CLK _12708_/D VGND VGND VPWR VPWR hold361/A sky130_fd_sc_hd__dfxtp_1
XFILLER_148_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13688_ _13700_/CLK _13688_/D repeater56/X VGND VGND VPWR VPWR _13688_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12639_ _14744_/Q _12637_/A _12638_/Y VGND VGND VPWR VPWR _14744_/D sky130_fd_sc_hd__o21a_1
XFILLER_157_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06160_ _06160_/A VGND VGND VPWR VPWR _14210_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold205 hold205/A VGND VGND VPWR VPWR hold205/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_14309_ _14543_/CLK _14309_/D VGND VGND VPWR VPWR _14309_/Q sky130_fd_sc_hd__dfxtp_1
X_06091_ _06091_/A VGND VGND VPWR VPWR _06105_/B sky130_fd_sc_hd__clkbuf_1
Xhold216 hold216/A VGND VGND VPWR VPWR hold216/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_160_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold227 hold227/A VGND VGND VPWR VPWR hold227/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold238 hold238/A VGND VGND VPWR VPWR hold238/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold249 hold249/A VGND VGND VPWR VPWR hold249/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09850_ _13683_/Q _13684_/Q VGND VGND VPWR VPWR _09858_/D sky130_fd_sc_hd__and2_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _13473_/D _08801_/B VGND VGND VPWR VPWR _11268_/B sky130_fd_sc_hd__xnor2_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06993_ _06990_/Y _06991_/X _06986_/A _06987_/Y VGND VGND VPWR VPWR _06993_/X sky130_fd_sc_hd__a211o_1
XFILLER_86_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09781_ _09781_/A VGND VGND VPWR VPWR _09781_/Y sky130_fd_sc_hd__inv_2
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05944_ _05944_/A _05944_/B _05944_/C VGND VGND VPWR VPWR _05945_/D sky130_fd_sc_hd__or3_1
X_08732_ _08724_/A _08728_/X _08741_/C VGND VGND VPWR VPWR _08739_/B sky130_fd_sc_hd__a21oi_1
XFILLER_26_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08663_ _08664_/A _08664_/B _08664_/C VGND VGND VPWR VPWR _08663_/X sky130_fd_sc_hd__a21o_1
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07614_ _07614_/A _07614_/B VGND VGND VPWR VPWR _07620_/B sky130_fd_sc_hd__xnor2_1
XFILLER_42_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08594_ _08544_/X _08671_/B _08671_/A VGND VGND VPWR VPWR _08596_/A sky130_fd_sc_hd__o21ai_2
XFILLER_81_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07545_ _09277_/B VGND VGND VPWR VPWR _09284_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_127_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _13963_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07476_ _07399_/X _07465_/Y _07475_/X VGND VGND VPWR VPWR _13147_/D sky130_fd_sc_hd__a21o_1
XFILLER_22_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09215_ _09215_/A VGND VGND VPWR VPWR _09215_/X sky130_fd_sc_hd__clkbuf_2
X_06427_ _06425_/X _06563_/C _06427_/S VGND VGND VPWR VPWR _06524_/C sky130_fd_sc_hd__mux2_1
XFILLER_22_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09146_ _13531_/Q _07365_/X _09161_/B VGND VGND VPWR VPWR _09146_/X sky130_fd_sc_hd__a21o_1
X_06358_ _14687_/Q _12874_/D VGND VGND VPWR VPWR _06358_/X sky130_fd_sc_hd__and2_1
XFILLER_148_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09077_ _09600_/A VGND VGND VPWR VPWR _09587_/S sky130_fd_sc_hd__clkbuf_4
X_06289_ _14186_/Q _14178_/Q _06289_/S VGND VGND VPWR VPWR _06289_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08028_ _12953_/Q _13253_/Q _10818_/B VGND VGND VPWR VPWR _08029_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09979_ _14429_/Q _14594_/Q _13754_/Q VGND VGND VPWR VPWR _09980_/B sky130_fd_sc_hd__mux2_1
XFILLER_103_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12990_ _14643_/CLK _12990_/D VGND VGND VPWR VPWR _13112_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_29_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11941_ _11941_/A VGND VGND VPWR VPWR _14276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _14716_/CLK _14660_/D VGND VGND VPWR VPWR _14660_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _11872_/A VGND VGND VPWR VPWR _14233_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13611_ _13622_/CLK _13611_/D repeater57/X VGND VGND VPWR VPWR _13611_/Q sky130_fd_sc_hd__dfrtp_2
X_10823_ _13131_/Q _10893_/A VGND VGND VPWR VPWR _10824_/A sky130_fd_sc_hd__and2_1
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14591_ _14644_/CLK _14591_/D VGND VGND VPWR VPWR _14591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_118_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _13653_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13542_ _13558_/CLK _13542_/D _12609_/A VGND VGND VPWR VPWR _13542_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_158_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10754_ _10754_/A VGND VGND VPWR VPWR _13041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10685_ _12879_/Q _10687_/B VGND VGND VPWR VPWR _10686_/A sky130_fd_sc_hd__and2_1
X_13473_ _14256_/CLK _13473_/D VGND VGND VPWR VPWR _13473_/Q sky130_fd_sc_hd__dfxtp_1
X_12424_ _12484_/A _12484_/B input6/X VGND VGND VPWR VPWR _12425_/A sky130_fd_sc_hd__and3_1
XFILLER_127_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12355_ _12377_/A VGND VGND VPWR VPWR _12364_/S sky130_fd_sc_hd__buf_2
XFILLER_142_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11306_ _11306_/A VGND VGND VPWR VPWR _13762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12286_ _12286_/A VGND VGND VPWR VPWR _14559_/D sky130_fd_sc_hd__clkbuf_1
X_11237_ _14617_/Q _14579_/Q _14510_/Q _14462_/Q _11186_/X _11187_/X VGND VGND VPWR
+ VPWR _11238_/A sky130_fd_sc_hd__mux4_1
XFILLER_4_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14025_ _14713_/CLK _14025_/D VGND VGND VPWR VPWR _14025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11168_ _11179_/A _11168_/B VGND VGND VPWR VPWR _11168_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10119_ _06152_/X _06289_/X _10119_/S VGND VGND VPWR VPWR _10120_/A sky130_fd_sc_hd__mux2_1
X_11099_ _14306_/Q _14476_/Q _14232_/Q _14062_/Q _11066_/X _11067_/X VGND VGND VPWR
+ VPWR _11099_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13809_ _13811_/CLK _13809_/D VGND VGND VPWR VPWR _13809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_109_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _13605_/CLK sky130_fd_sc_hd__clkbuf_16
X_07330_ _07428_/A _07328_/X _07329_/Y VGND VGND VPWR VPWR _07330_/X sky130_fd_sc_hd__o21ba_1
XFILLER_32_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07261_ _08157_/A _07261_/B _09086_/C VGND VGND VPWR VPWR _07261_/X sky130_fd_sc_hd__and3_1
X_09000_ _08995_/A _08994_/B _08996_/B _08996_/A VGND VGND VPWR VPWR _09003_/A sky130_fd_sc_hd__a22o_1
X_06212_ hold94/A VGND VGND VPWR VPWR _06321_/S sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_7_0_clk clkbuf_3_7_0_clk/A VGND VGND VPWR VPWR clkbuf_3_7_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07192_ _07204_/A _07204_/B VGND VGND VPWR VPWR _07201_/A sky130_fd_sc_hd__xnor2_1
X_06143_ _14190_/Q _14182_/Q _06289_/S VGND VGND VPWR VPWR _06146_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06074_ hold498/A _06075_/C _06075_/D _06076_/A VGND VGND VPWR VPWR _06259_/B sky130_fd_sc_hd__and4_1
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09902_ _09902_/A VGND VGND VPWR VPWR _13698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09833_ _09840_/A _09833_/B VGND VGND VPWR VPWR _09833_/Y sky130_fd_sc_hd__xnor2_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _09760_/B _09763_/Y _09774_/S VGND VGND VPWR VPWR _09765_/A sky130_fd_sc_hd__mux2_1
X_06976_ _06976_/A VGND VGND VPWR VPWR _06976_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_55_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08715_ _08742_/A VGND VGND VPWR VPWR _08715_/Y sky130_fd_sc_hd__inv_2
X_05927_ _13720_/Q _13729_/Q _13730_/Q _13731_/Q VGND VGND VPWR VPWR _05928_/C sky130_fd_sc_hd__and4_1
XFILLER_100_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09695_ _13669_/Q _09695_/B VGND VGND VPWR VPWR _09696_/B sky130_fd_sc_hd__nand2_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08646_ _08546_/Y _08645_/Y _08544_/X VGND VGND VPWR VPWR _08646_/Y sky130_fd_sc_hd__o21ai_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08577_ _13443_/Q _08577_/B VGND VGND VPWR VPWR _08590_/A sky130_fd_sc_hd__nand2_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07528_ _13154_/Q _09237_/B VGND VGND VPWR VPWR _07530_/C sky130_fd_sc_hd__xor2_1
XFILLER_22_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07459_ _07457_/Y _07443_/B _07454_/C _07458_/Y _07452_/B VGND VGND VPWR VPWR _07459_/X
+ sky130_fd_sc_hd__o32a_1
X_10470_ _10438_/B _10462_/A _10452_/A _10452_/B VGND VGND VPWR VPWR _10471_/B sky130_fd_sc_hd__o22ai_2
XFILLER_6_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09129_ _09125_/X _09128_/Y _07359_/X VGND VGND VPWR VPWR _13530_/D sky130_fd_sc_hd__a21o_1
XFILLER_109_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12140_ _12140_/A VGND VGND VPWR VPWR _14484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12071_ _12071_/A VGND VGND VPWR VPWR _14453_/D sky130_fd_sc_hd__clkbuf_1
X_11022_ _14262_/Q _14653_/Q _13760_/Q _14708_/Q _11020_/X _11021_/X VGND VGND VPWR
+ VPWR _11023_/B sky130_fd_sc_hd__mux4_1
XFILLER_77_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12973_ _12974_/CLK hold170/X VGND VGND VPWR VPWR _12973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14712_ _14712_/CLK _14712_/D VGND VGND VPWR VPWR _14712_/Q sky130_fd_sc_hd__dfxtp_1
X_11924_ _11924_/A VGND VGND VPWR VPWR _14268_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _14643_/CLK _14643_/D VGND VGND VPWR VPWR _14643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _11877_/A VGND VGND VPWR VPWR _11864_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10806_ _13023_/Q _10812_/B VGND VGND VPWR VPWR _10807_/A sky130_fd_sc_hd__and2_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14574_ _14733_/CLK _14574_/D VGND VGND VPWR VPWR _14574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11786_ _11834_/B VGND VGND VPWR VPWR _11795_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_13_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13525_ _13525_/CLK _13525_/D _12609_/A VGND VGND VPWR VPWR _13525_/Q sky130_fd_sc_hd__dfrtp_1
X_10737_ _10737_/A VGND VGND VPWR VPWR _12945_/D sky130_fd_sc_hd__clkbuf_1
X_13456_ _13605_/CLK _13456_/D repeater57/X VGND VGND VPWR VPWR _13456_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_127_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10668_ _10671_/C _10668_/B VGND VGND VPWR VPWR _12915_/D sky130_fd_sc_hd__nor2_1
X_12407_ _12502_/A VGND VGND VPWR VPWR _12418_/A sky130_fd_sc_hd__clkbuf_1
X_10599_ _14639_/Q _12336_/C _14640_/Q _14646_/Q VGND VGND VPWR VPWR _10600_/A sky130_fd_sc_hd__or4b_1
X_13387_ _13423_/CLK _13387_/D VGND VGND VPWR VPWR _13387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12338_ _14641_/Q _12340_/B VGND VGND VPWR VPWR _12339_/A sky130_fd_sc_hd__and2_1
XFILLER_154_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14762__73 VGND VGND VPWR VPWR _14762__73/HI _13033_/D sky130_fd_sc_hd__conb_1
XFILLER_99_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12269_ _12269_/A VGND VGND VPWR VPWR _14549_/D sky130_fd_sc_hd__clkbuf_1
X_14008_ _14012_/CLK _14008_/D VGND VGND VPWR VPWR _14008_/Q sky130_fd_sc_hd__dfxtp_1
X_06830_ _06796_/A _06800_/B _06813_/C _06769_/B VGND VGND VPWR VPWR _06840_/A sky130_fd_sc_hd__o31a_2
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06761_ _06775_/A _06740_/X VGND VGND VPWR VPWR _06762_/B sky130_fd_sc_hd__or2b_1
XFILLER_48_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08500_ _08500_/A _08500_/B VGND VGND VPWR VPWR _08500_/X sky130_fd_sc_hd__xor2_1
XFILLER_64_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09480_ _13604_/Q _09472_/B _09478_/B _09479_/Y VGND VGND VPWR VPWR _09480_/Y sky130_fd_sc_hd__a22oi_1
X_06692_ _07804_/B _06690_/B _06689_/X VGND VGND VPWR VPWR _06696_/B sky130_fd_sc_hd__o21bai_1
XFILLER_63_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08431_ _13471_/Q _13476_/Q VGND VGND VPWR VPWR _08431_/X sky130_fd_sc_hd__and2b_1
XFILLER_24_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08362_ _13079_/Q _13360_/Q _08362_/S VGND VGND VPWR VPWR _08363_/A sky130_fd_sc_hd__mux2_1
X_07313_ _07313_/A _07335_/A VGND VGND VPWR VPWR _09112_/B sky130_fd_sc_hd__and2_1
X_08293_ _13370_/Q _13371_/Q VGND VGND VPWR VPWR _08301_/D sky130_fd_sc_hd__and2_1
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07244_ _13658_/Q _13656_/Q _07299_/S VGND VGND VPWR VPWR _07244_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07175_ _07149_/A _07175_/B VGND VGND VPWR VPWR _07175_/X sky130_fd_sc_hd__and2b_1
XFILLER_117_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06126_ _14203_/Q _14201_/Q _10107_/A VGND VGND VPWR VPWR _06126_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06057_ _06057_/A VGND VGND VPWR VPWR _10019_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09816_ _09816_/A _09816_/B VGND VGND VPWR VPWR _09816_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09747_ _13673_/Q _09748_/B VGND VGND VPWR VPWR _09749_/A sky130_fd_sc_hd__and2_1
XFILLER_36_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06959_ _13023_/Q _07981_/B VGND VGND VPWR VPWR _06967_/B sky130_fd_sc_hd__xor2_1
XFILLER_27_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _09720_/A _13667_/Q _09678_/C VGND VGND VPWR VPWR _09682_/A sky130_fd_sc_hd__and3_1
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08629_ _08630_/B _08630_/C _08630_/D _08630_/A VGND VGND VPWR VPWR _08629_/X sky130_fd_sc_hd__a31o_1
XFILLER_54_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11640_/A VGND VGND VPWR VPWR _13995_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11571_ _11571_/A VGND VGND VPWR VPWR _13867_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13310_ _14275_/CLK hold368/X VGND VGND VPWR VPWR _13310_/Q sky130_fd_sc_hd__dfxtp_1
X_10522_ _12990_/D VGND VGND VPWR VPWR _10557_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14290_ _14292_/CLK _14290_/D VGND VGND VPWR VPWR hold283/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10453_ _10453_/A _10453_/B VGND VGND VPWR VPWR _14007_/D sky130_fd_sc_hd__xnor2_1
XFILLER_108_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13241_ _14010_/CLK _13241_/D VGND VGND VPWR VPWR _13513_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_136_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10384_ _13518_/Q _10393_/A VGND VGND VPWR VPWR _10405_/A sky130_fd_sc_hd__and2_1
XFILLER_151_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13172_ _13524_/CLK _13172_/D VGND VGND VPWR VPWR _13172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12123_ _12123_/A VGND VGND VPWR VPWR _14476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12054_ _12076_/A VGND VGND VPWR VPWR _12063_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_77_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11005_ _11037_/A _11005_/B VGND VGND VPWR VPWR _11005_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12956_ _13039_/CLK hold423/X VGND VGND VPWR VPWR _12956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11907_ _14261_/Q _11462_/X _11907_/S VGND VGND VPWR VPWR _11908_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _12930_/CLK _12887_/D hold1/X VGND VGND VPWR VPWR _12887_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _14647_/CLK _14626_/D VGND VGND VPWR VPWR _14626_/Q sky130_fd_sc_hd__dfxtp_1
X_11838_ _14148_/D _14149_/D _14151_/D _14153_/D VGND VGND VPWR VPWR _11839_/C sky130_fd_sc_hd__or4_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _14557_/CLK _14557_/D VGND VGND VPWR VPWR _14557_/Q sky130_fd_sc_hd__dfxtp_1
X_11769_ _11769_/A VGND VGND VPWR VPWR _14079_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_40_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _13258_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_146_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13508_ _13698_/CLK hold263/X VGND VGND VPWR VPWR _13508_/Q sky130_fd_sc_hd__dfxtp_1
X_14488_ _14726_/CLK _14488_/D VGND VGND VPWR VPWR _14488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13439_ _13598_/CLK _13439_/D repeater56/X VGND VGND VPWR VPWR _13439_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_127_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08980_ _08992_/A _08992_/B VGND VGND VPWR VPWR _08989_/A sky130_fd_sc_hd__xnor2_1
XFILLER_130_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07931_ _07934_/A _07949_/B VGND VGND VPWR VPWR _07931_/X sky130_fd_sc_hd__xor2_1
XFILLER_69_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07862_ _07862_/A VGND VGND VPWR VPWR _13260_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09601_ _13398_/Q _13596_/Q _09609_/S VGND VGND VPWR VPWR _09602_/A sky130_fd_sc_hd__mux2_2
X_06813_ _06813_/A _06813_/B _06813_/C VGND VGND VPWR VPWR _06881_/C sky130_fd_sc_hd__or3_1
XFILLER_113_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07793_ _07793_/A VGND VGND VPWR VPWR _13664_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09532_ _09532_/A _09532_/B _09532_/C VGND VGND VPWR VPWR _09532_/X sky130_fd_sc_hd__or3_1
X_06744_ _06703_/X _07856_/B _06740_/X _06743_/Y VGND VGND VPWR VPWR _13004_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09463_ _13603_/Q _09464_/B VGND VGND VPWR VPWR _09475_/A sky130_fd_sc_hd__nand2_1
X_06675_ _06852_/A _06672_/X _06674_/X VGND VGND VPWR VPWR _06675_/X sky130_fd_sc_hd__a21o_1
XFILLER_51_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08414_ _13102_/Q _13383_/Q _08418_/S VGND VGND VPWR VPWR _08415_/A sky130_fd_sc_hd__mux2_1
X_09394_ _13593_/Q _09394_/B VGND VGND VPWR VPWR _09396_/A sky130_fd_sc_hd__nand2_2
XFILLER_149_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08345_ _13385_/Q _08340_/X _08344_/Y VGND VGND VPWR VPWR _13385_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_31_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _13031_/CLK sky130_fd_sc_hd__clkbuf_16
X_08276_ _08283_/A _08276_/B VGND VGND VPWR VPWR _08276_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_137_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07227_ _13657_/Q _13655_/Q _07299_/S VGND VGND VPWR VPWR _07227_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07158_ _07158_/A VGND VGND VPWR VPWR _13348_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06109_ _13787_/Q _13788_/Q _13789_/Q _13790_/Q VGND VGND VPWR VPWR _06109_/X sky130_fd_sc_hd__or4_1
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07089_ _07119_/B _07141_/B hold154/A _07119_/A VGND VGND VPWR VPWR _07093_/A sky130_fd_sc_hd__a22oi_2
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_98_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _13727_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_120_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12810_ _13622_/CLK _12810_/D VGND VGND VPWR VPWR hold100/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13790_ _13799_/CLK _13790_/D VGND VGND VPWR VPWR _13790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _13423_/CLK _12741_/D VGND VGND VPWR VPWR hold477/A sky130_fd_sc_hd__dfxtp_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _13353_/CLK _12672_/D VGND VGND VPWR VPWR _12672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _14413_/CLK hold94/X VGND VGND VPWR VPWR _14411_/Q sky130_fd_sc_hd__dfxtp_1
X_11623_ _13988_/Q _11478_/X _11623_/S VGND VGND VPWR VPWR _11624_/A sky130_fd_sc_hd__mux2_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_22_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _13554_/CLK sky130_fd_sc_hd__clkbuf_16
X_14342_ _14697_/CLK hold482/X VGND VGND VPWR VPWR _14342_/Q sky130_fd_sc_hd__dfxtp_1
X_11554_ _11576_/A VGND VGND VPWR VPWR _11563_/B sky130_fd_sc_hd__clkbuf_1
X_10505_ _10438_/B _10439_/A _10504_/Y VGND VGND VPWR VPWR _14005_/D sky130_fd_sc_hd__a21oi_1
XFILLER_7_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14273_ _14720_/CLK _14273_/D VGND VGND VPWR VPWR _14273_/Q sky130_fd_sc_hd__dfxtp_1
X_11485_ _14516_/Q VGND VGND VPWR VPWR _11485_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13224_ _13606_/CLK hold471/X VGND VGND VPWR VPWR _13224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10436_ hold46/A VGND VGND VPWR VPWR _10441_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13155_ _14530_/CLK _13155_/D _12609_/A VGND VGND VPWR VPWR _13155_/Q sky130_fd_sc_hd__dfrtp_2
X_10367_ _10367_/A VGND VGND VPWR VPWR _14213_/D sky130_fd_sc_hd__clkbuf_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _14469_/Q _11965_/X _12106_/S VGND VGND VPWR VPWR _12107_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10298_ _14681_/Q _14682_/Q _14688_/Q _12030_/C VGND VGND VPWR VPWR _10299_/A sky130_fd_sc_hd__or4_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ _13565_/CLK hold417/X VGND VGND VPWR VPWR _13086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_89_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _14212_/CLK sky130_fd_sc_hd__clkbuf_16
X_12037_ _12037_/A VGND VGND VPWR VPWR _14383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13988_ _14709_/CLK _13988_/D VGND VGND VPWR VPWR _13988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12939_ _12974_/CLK _12939_/D VGND VGND VPWR VPWR hold194/A sky130_fd_sc_hd__dfxtp_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06460_ _06471_/A _06460_/B _06460_/C VGND VGND VPWR VPWR _06462_/B sky130_fd_sc_hd__and3_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14609_ _14610_/CLK _14609_/D VGND VGND VPWR VPWR _14609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06391_ _06391_/A _06391_/B VGND VGND VPWR VPWR _12876_/D sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_13_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _14319_/CLK sky130_fd_sc_hd__clkbuf_16
X_08130_ _13425_/Q VGND VGND VPWR VPWR _08228_/S sky130_fd_sc_hd__inv_2
XFILLER_159_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08061_ _08061_/A VGND VGND VPWR VPWR _12691_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07012_ _07040_/A _07031_/A VGND VGND VPWR VPWR _07013_/B sky130_fd_sc_hd__nand2_1
XFILLER_146_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08963_ _08937_/A _08963_/B VGND VGND VPWR VPWR _08963_/X sky130_fd_sc_hd__and2b_1
XFILLER_88_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07914_ _07914_/A _07914_/B _07916_/B VGND VGND VPWR VPWR _07914_/Y sky130_fd_sc_hd__nand3_1
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08894_ _08894_/A _08894_/B VGND VGND VPWR VPWR _08911_/A sky130_fd_sc_hd__nand2_1
XFILLER_111_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07845_ _07846_/B _07846_/C _13259_/Q VGND VGND VPWR VPWR _07847_/A sky130_fd_sc_hd__a21oi_1
X_07776_ _07783_/A _07776_/B VGND VGND VPWR VPWR _07778_/C sky130_fd_sc_hd__xnor2_1
XFILLER_71_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09515_ _09534_/A _09508_/Y _09510_/X _08542_/A VGND VGND VPWR VPWR _09515_/Y sky130_fd_sc_hd__a31oi_1
X_06727_ _06727_/A _06727_/B VGND VGND VPWR VPWR _06731_/A sky130_fd_sc_hd__or2_1
XFILLER_52_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09446_ _09447_/D _09454_/B _09446_/C _09454_/D VGND VGND VPWR VPWR _09446_/X sky130_fd_sc_hd__or4_1
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06658_ _07804_/B _07804_/C _12999_/Q VGND VGND VPWR VPWR _06659_/B sky130_fd_sc_hd__a21oi_1
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09377_ _09377_/A _09377_/B _09377_/C VGND VGND VPWR VPWR _09377_/Y sky130_fd_sc_hd__nand3_1
X_06589_ _12896_/Q _06595_/B _06542_/X VGND VGND VPWR VPWR _06590_/B sky130_fd_sc_hd__o21ai_1
X_08328_ _08331_/B _09084_/A _08328_/C VGND VGND VPWR VPWR _08329_/A sky130_fd_sc_hd__and3b_1
XFILLER_153_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08259_ _08259_/A VGND VGND VPWR VPWR _13366_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11270_ _10635_/B _11270_/B VGND VGND VPWR VPWR _11271_/A sky130_fd_sc_hd__and2b_1
XFILLER_4_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10221_ _10221_/A VGND VGND VPWR VPWR _14398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10152_ _14287_/D _10151_/X _10179_/S VGND VGND VPWR VPWR _10153_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10083_ _10078_/X _10082_/X _14048_/D VGND VGND VPWR VPWR _10084_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_13911_ _13978_/CLK _13911_/D VGND VGND VPWR VPWR _13911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13842_ _14724_/CLK _13842_/D VGND VGND VPWR VPWR _13842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13773_ _14721_/CLK _13773_/D VGND VGND VPWR VPWR _13773_/Q sky130_fd_sc_hd__dfxtp_1
X_10985_ _10985_/A VGND VGND VPWR VPWR _10985_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12724_ _13606_/CLK _12724_/D VGND VGND VPWR VPWR hold485/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12655_ _14082_/CLK hold501/X _12609_/A VGND VGND VPWR VPWR hold512/A sky130_fd_sc_hd__dfrtp_1
XFILLER_90_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11606_ _13980_/Q _11453_/X _11612_/S VGND VGND VPWR VPWR _11607_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12586_ _12586_/A _14730_/Q VGND VGND VPWR VPWR _12586_/Y sky130_fd_sc_hd__nand2_1
X_14325_ _14688_/CLK _14325_/D VGND VGND VPWR VPWR _14325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11537_ _13628_/Q _11541_/B VGND VGND VPWR VPWR _11538_/A sky130_fd_sc_hd__and2_1
XFILLER_144_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold409 hold409/A VGND VGND VPWR VPWR hold409/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_109_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14256_ _14256_/CLK _14256_/D VGND VGND VPWR VPWR _14256_/Q sky130_fd_sc_hd__dfxtp_1
X_11468_ _11468_/A VGND VGND VPWR VPWR _13824_/D sky130_fd_sc_hd__clkbuf_1
X_13207_ _14012_/CLK hold360/X VGND VGND VPWR VPWR _13207_/Q sky130_fd_sc_hd__dfxtp_1
X_10419_ _10426_/A _10419_/B VGND VGND VPWR VPWR _10421_/C sky130_fd_sc_hd__nor2_1
X_14187_ _14201_/CLK _14187_/D VGND VGND VPWR VPWR _14187_/Q sky130_fd_sc_hd__dfxtp_1
X_11399_ _13723_/Q _11405_/B VGND VGND VPWR VPWR _11400_/A sky130_fd_sc_hd__and2_1
XFILLER_98_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _13434_/CLK _13138_/D repeater56/X VGND VGND VPWR VPWR _13138_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05960_ _13631_/Q _13632_/Q _13633_/Q _13634_/Q VGND VGND VPWR VPWR _05963_/C sky130_fd_sc_hd__or4_1
X_13069_ _14082_/CLK _13069_/D VGND VGND VPWR VPWR hold250/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_2_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _14615_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07630_ _07641_/B _07656_/B VGND VGND VPWR VPWR _07631_/B sky130_fd_sc_hd__nor2_1
XFILLER_93_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07561_ _09250_/B VGND VGND VPWR VPWR _09271_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09300_ _09300_/A VGND VGND VPWR VPWR _12778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06512_ _06554_/C VGND VGND VPWR VPWR _06563_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07492_ _07493_/A _07493_/B _07504_/C VGND VGND VPWR VPWR _07498_/B sky130_fd_sc_hd__a21o_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09231_ _09125_/X _09230_/Y _07475_/X VGND VGND VPWR VPWR _13544_/D sky130_fd_sc_hd__a21o_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06443_ _13107_/D _06444_/A VGND VGND VPWR VPWR _06443_/X sky130_fd_sc_hd__or2b_1
XFILLER_159_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09162_ _09135_/A _09135_/B _09135_/C _09161_/X _09160_/B VGND VGND VPWR VPWR _09162_/X
+ sky130_fd_sc_hd__a311o_1
X_06374_ hold41/X _13389_/D _06373_/X VGND VGND VPWR VPWR _14647_/D sky130_fd_sc_hd__o21ba_1
XFILLER_148_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08113_ _08113_/A _08113_/B VGND VGND VPWR VPWR _13354_/D sky130_fd_sc_hd__xor2_1
X_09093_ _13525_/Q _09093_/B VGND VGND VPWR VPWR _09095_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08044_ _08044_/A VGND VGND VPWR VPWR _12683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09995_ _10636_/A _14625_/Q VGND VGND VPWR VPWR _11270_/B sky130_fd_sc_hd__and2b_1
XFILLER_142_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08946_ _08946_/A VGND VGND VPWR VPWR _14251_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08877_ _08907_/B _08929_/B _13431_/Q _08907_/A VGND VGND VPWR VPWR _08881_/A sky130_fd_sc_hd__a22oi_2
XFILLER_57_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07828_ _07833_/A _07828_/B VGND VGND VPWR VPWR _07829_/B sky130_fd_sc_hd__and2b_1
XFILLER_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07759_ _07760_/A _07760_/B _07759_/C VGND VGND VPWR VPWR _07778_/A sky130_fd_sc_hd__or3_1
XFILLER_53_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10770_ _10781_/A VGND VGND VPWR VPWR _10779_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09429_ _09447_/C _09454_/A _09427_/X _09365_/A VGND VGND VPWR VPWR _09429_/X sky130_fd_sc_hd__o31a_1
XFILLER_9_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12440_ _12440_/A VGND VGND VPWR VPWR _14652_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12371_ _14608_/Q _11991_/X _12375_/S VGND VGND VPWR VPWR _12372_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14110_ _14209_/CLK hold87/X VGND VGND VPWR VPWR _14110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11322_ _11322_/A VGND VGND VPWR VPWR _13767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14041_ _14050_/CLK _14041_/D VGND VGND VPWR VPWR _14041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11253_ _12626_/B _11253_/B VGND VGND VPWR VPWR _11253_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10204_ _10626_/D _10203_/X _10206_/S VGND VGND VPWR VPWR _10205_/A sky130_fd_sc_hd__mux2_1
X_11184_ _11136_/X _11181_/X _11183_/X _11157_/X VGND VGND VPWR VPWR _11184_/X sky130_fd_sc_hd__o211a_1
XFILLER_106_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10135_ _13868_/Q _13852_/Q _10137_/S VGND VGND VPWR VPWR _10136_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10066_ _10066_/A VGND VGND VPWR VPWR _14046_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13825_ _14737_/CLK _13825_/D VGND VGND VPWR VPWR _13825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13756_ _14704_/CLK _13756_/D VGND VGND VPWR VPWR _13756_/Q sky130_fd_sc_hd__dfxtp_1
X_10968_ _12649_/B VGND VGND VPWR VPWR _11037_/A sky130_fd_sc_hd__buf_2
XFILLER_43_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12707_ _14098_/CLK _12707_/D VGND VGND VPWR VPWR hold332/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13687_ _13700_/CLK _13687_/D repeater56/X VGND VGND VPWR VPWR _13687_/Q sky130_fd_sc_hd__dfrtp_1
X_10899_ _10899_/A _10899_/B _10899_/C _10899_/D VGND VGND VPWR VPWR _10901_/A sky130_fd_sc_hd__or4_1
X_12638_ _14744_/Q _12637_/A _12633_/B VGND VGND VPWR VPWR _12638_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_129_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12569_ _14743_/Q VGND VGND VPWR VPWR _12569_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14308_ _14543_/CLK _14308_/D VGND VGND VPWR VPWR _14308_/Q sky130_fd_sc_hd__dfxtp_1
X_06090_ _06090_/A VGND VGND VPWR VPWR _13978_/D sky130_fd_sc_hd__clkbuf_1
Xhold206 hold206/A VGND VGND VPWR VPWR hold206/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold217 hold217/A VGND VGND VPWR VPWR hold217/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold228 hold228/A VGND VGND VPWR VPWR hold228/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_160_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14239_ _14510_/CLK _14239_/D VGND VGND VPWR VPWR _14239_/Q sky130_fd_sc_hd__dfxtp_1
Xhold239 hold239/A VGND VGND VPWR VPWR hold239/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _08828_/A _08819_/A VGND VGND VPWR VPWR _08801_/B sky130_fd_sc_hd__nand2_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09780_ _09780_/A _09793_/A VGND VGND VPWR VPWR _09783_/A sky130_fd_sc_hd__or2_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06992_ _06986_/A _06987_/Y _06990_/Y _06991_/X VGND VGND VPWR VPWR _06992_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_112_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _08739_/A _08731_/B VGND VGND VPWR VPWR _08741_/C sky130_fd_sc_hd__or2_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05943_ _13867_/Q _13868_/Q _13869_/Q _13870_/Q VGND VGND VPWR VPWR _05944_/C sky130_fd_sc_hd__or4_1
XFILLER_100_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08662_ _08662_/A _08662_/B VGND VGND VPWR VPWR _08664_/C sky130_fd_sc_hd__or2_2
XFILLER_53_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07613_ _07613_/A _07723_/A VGND VGND VPWR VPWR _07614_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08593_ _08589_/Y _08590_/X _08592_/X _08517_/X VGND VGND VPWR VPWR _13444_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07544_ _07399_/X _07543_/X _07475_/X VGND VGND VPWR VPWR _13156_/D sky130_fd_sc_hd__a21o_1
XFILLER_34_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07475_ _07499_/A VGND VGND VPWR VPWR _07475_/X sky130_fd_sc_hd__buf_2
XFILLER_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09214_ _09214_/A _09214_/B _09220_/D VGND VGND VPWR VPWR _09214_/Y sky130_fd_sc_hd__nand3_1
XFILLER_10_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06426_ _06469_/A _12671_/Q VGND VGND VPWR VPWR _06563_/C sky130_fd_sc_hd__and2_1
XFILLER_148_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09145_ _13533_/Q _09151_/B VGND VGND VPWR VPWR _09159_/A sky130_fd_sc_hd__xnor2_1
X_06357_ _14687_/Q _12874_/D VGND VGND VPWR VPWR _06357_/Y sky130_fd_sc_hd__nor2_1
XFILLER_136_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06288_ _13953_/D _13956_/D _06284_/X hold503/X VGND VGND VPWR VPWR _13961_/D sky130_fd_sc_hd__o31ai_1
X_09076_ _09076_/A VGND VGND VPWR VPWR _12771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08027_ _08027_/A VGND VGND VPWR VPWR _12673_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09978_ _10597_/A _14591_/Q VGND VGND VPWR VPWR _12404_/B sky130_fd_sc_hd__and2b_1
XFILLER_58_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08929_ _08929_/A _08929_/B _08929_/C _08951_/B VGND VGND VPWR VPWR _08930_/B sky130_fd_sc_hd__and4_1
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11940_ _14276_/Q _11510_/X _11940_/S VGND VGND VPWR VPWR _11941_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _14233_/Q _11488_/X _11875_/S VGND VGND VPWR VPWR _11872_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _13610_/CLK _13610_/D repeater57/X VGND VGND VPWR VPWR _13610_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10822_ _10822_/A VGND VGND VPWR VPWR _10893_/A sky130_fd_sc_hd__buf_2
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _14688_/CLK _14590_/D VGND VGND VPWR VPWR _14590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13541_ _13558_/CLK _13541_/D _12609_/A VGND VGND VPWR VPWR _13541_/Q sky130_fd_sc_hd__dfrtp_1
X_10753_ _12999_/Q _10820_/A VGND VGND VPWR VPWR _10754_/A sky130_fd_sc_hd__and2_1
XFILLER_41_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13472_ _13621_/CLK _13472_/D VGND VGND VPWR VPWR _13472_/Q sky130_fd_sc_hd__dfxtp_1
X_10684_ _10684_/A VGND VGND VPWR VPWR _12921_/D sky130_fd_sc_hd__clkbuf_1
X_12423_ _12423_/A VGND VGND VPWR VPWR _14644_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12354_ _12354_/A VGND VGND VPWR VPWR _14600_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11305_ _13762_/Q _11304_/X _11311_/S VGND VGND VPWR VPWR _11306_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12285_ _14559_/Q _11956_/X _12291_/S VGND VGND VPWR VPWR _12286_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14024_ _14713_/CLK _14024_/D VGND VGND VPWR VPWR _14024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11236_ _11207_/X _11233_/X _11235_/X _12647_/A VGND VGND VPWR VPWR _11236_/X sky130_fd_sc_hd__o211a_1
XFILLER_4_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11167_ _11159_/X _11161_/Y _11165_/Y _11166_/X VGND VGND VPWR VPWR _11168_/B sky130_fd_sc_hd__a211o_1
XFILLER_1_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10118_ _10118_/A VGND VGND VPWR VPWR _14201_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11098_ _13328_/Q _11079_/X _11087_/X _11097_/Y VGND VGND VPWR VPWR _13328_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10049_ _10049_/A VGND VGND VPWR VPWR _13950_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13808_ _13811_/CLK _13808_/D VGND VGND VPWR VPWR _13808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13739_ _13811_/CLK hold346/X VGND VGND VPWR VPWR _13739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07260_ _07473_/A VGND VGND VPWR VPWR _08157_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06211_ _14406_/Q _14398_/Q hold94/A VGND VGND VPWR VPWR _06215_/D sky130_fd_sc_hd__mux2_1
X_07191_ _07191_/A _07191_/B VGND VGND VPWR VPWR _07204_/B sky130_fd_sc_hd__nor2_1
X_06142_ _14194_/D VGND VGND VPWR VPWR _06289_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_118_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06073_ _13958_/Q _13950_/Q _06256_/S VGND VGND VPWR VPWR _06076_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09901_ _09899_/X _09901_/B VGND VGND VPWR VPWR _09902_/A sky130_fd_sc_hd__and2b_1
XFILLER_113_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ _09815_/A _09816_/A _09815_/B _09824_/A _09831_/X VGND VGND VPWR VPWR _09833_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _09763_/A _09763_/B VGND VGND VPWR VPWR _09763_/Y sky130_fd_sc_hd__xnor2_1
X_06975_ _06945_/X _06978_/B _06973_/Y _06974_/X VGND VGND VPWR VPWR _13024_/D sky130_fd_sc_hd__a31o_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08714_ _08714_/A _08714_/B _08714_/C _08714_/D VGND VGND VPWR VPWR _08742_/A sky130_fd_sc_hd__or4_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05926_ _13732_/Q _13737_/Q _13738_/Q _13739_/Q VGND VGND VPWR VPWR _05928_/B sky130_fd_sc_hd__and4_1
X_09694_ _13669_/Q _09695_/B VGND VGND VPWR VPWR _09696_/A sky130_fd_sc_hd__or2_1
XFILLER_66_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _08645_/A _08645_/B VGND VGND VPWR VPWR _08645_/Y sky130_fd_sc_hd__nor2_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08576_ _08517_/X _08577_/B _08590_/B _08575_/Y VGND VGND VPWR VPWR _13443_/D sky130_fd_sc_hd__a22o_1
XFILLER_70_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07527_ _07530_/B _07525_/X _07526_/X VGND VGND VPWR VPWR _13153_/D sky130_fd_sc_hd__o21bai_1
XFILLER_22_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07458_ _13145_/Q _09183_/B _07452_/A VGND VGND VPWR VPWR _07458_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_10_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06409_ _06444_/A VGND VGND VPWR VPWR _06482_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07389_ _07389_/A _07389_/B VGND VGND VPWR VPWR _07401_/B sky130_fd_sc_hd__or2_2
X_09128_ _09134_/D _09128_/B VGND VGND VPWR VPWR _09128_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09059_ _09059_/A VGND VGND VPWR VPWR _12763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12070_ _11320_/X _14453_/Q _12074_/S VGND VGND VPWR VPWR _12071_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11021_ _11092_/A VGND VGND VPWR VPWR _11021_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12972_ _12974_/CLK hold194/X VGND VGND VPWR VPWR _12972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11923_ _14268_/Q _11485_/X _11929_/S VGND VGND VPWR VPWR _11924_/A sky130_fd_sc_hd__mux2_1
X_14711_ _14712_/CLK _14711_/D VGND VGND VPWR VPWR _14711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _14643_/CLK _14642_/D VGND VGND VPWR VPWR _14642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ _11854_/A VGND VGND VPWR VPWR _14225_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _10805_/A VGND VGND VPWR VPWR _13064_/D sky130_fd_sc_hd__clkbuf_1
X_14573_ _14619_/CLK _14573_/D VGND VGND VPWR VPWR _14573_/Q sky130_fd_sc_hd__dfxtp_1
X_11785_ _11785_/A VGND VGND VPWR VPWR _14086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13524_ _13524_/CLK _13524_/D hold1/X VGND VGND VPWR VPWR _13524_/Q sky130_fd_sc_hd__dfrtp_1
X_10736_ _12902_/Q _10742_/B VGND VGND VPWR VPWR _10737_/A sky130_fd_sc_hd__and2_1
X_13455_ _13700_/CLK _13455_/D repeater57/X VGND VGND VPWR VPWR _13455_/Q sky130_fd_sc_hd__dfrtp_1
X_10667_ _14340_/Q _10665_/A _10656_/X VGND VGND VPWR VPWR _10668_/B sky130_fd_sc_hd__o21ai_1
X_12406_ input28/X VGND VGND VPWR VPWR _12502_/A sky130_fd_sc_hd__buf_2
XFILLER_139_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13386_ _13423_/CLK _13386_/D repeater56/X VGND VGND VPWR VPWR _13386_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10598_ _14629_/Q _14633_/Q VGND VGND VPWR VPWR _14623_/D sky130_fd_sc_hd__xor2_1
X_12337_ _12337_/A VGND VGND VPWR VPWR _14592_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12268_ _11348_/X _14549_/Q _12270_/S VGND VGND VPWR VPWR _12269_/A sky130_fd_sc_hd__mux2_1
X_14007_ _14679_/CLK _14007_/D VGND VGND VPWR VPWR _14007_/Q sky130_fd_sc_hd__dfxtp_1
X_11219_ _11242_/A _11219_/B VGND VGND VPWR VPWR _11219_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12199_ _12199_/A VGND VGND VPWR VPWR _14510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06760_ _13004_/Q _07856_/B VGND VGND VPWR VPWR _06775_/A sky130_fd_sc_hd__and2_1
XFILLER_48_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06691_ _06786_/A VGND VGND VPWR VPWR _06719_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08430_ _14247_/Q _14245_/Q _08506_/S VGND VGND VPWR VPWR _08430_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08361_ _08361_/A VGND VGND VPWR VPWR _12714_/D sky130_fd_sc_hd__clkbuf_1
X_07312_ _07350_/A _07349_/A VGND VGND VPWR VPWR _07335_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08292_ _13370_/Q _08294_/A _08291_/Y VGND VGND VPWR VPWR _13370_/D sky130_fd_sc_hd__o21a_1
X_07243_ _13662_/Q _13660_/Q _13170_/Q VGND VGND VPWR VPWR _07243_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07174_ _07174_/A _07174_/B VGND VGND VPWR VPWR _07178_/B sky130_fd_sc_hd__and2_1
XFILLER_145_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06125_ _14209_/Q VGND VGND VPWR VPWR _10107_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06056_ _13971_/Q _13969_/Q _10020_/A VGND VGND VPWR VPWR _06056_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09815_ _09815_/A _09815_/B VGND VGND VPWR VPWR _09816_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09746_ _09758_/A _09746_/B _09746_/C VGND VGND VPWR VPWR _09748_/B sky130_fd_sc_hd__and3_1
XFILLER_39_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06958_ _06956_/Y _06957_/X _06897_/X VGND VGND VPWR VPWR _13022_/D sky130_fd_sc_hd__a21o_1
XFILLER_100_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05909_ _05909_/A _05909_/B _05909_/C VGND VGND VPWR VPWR _05910_/D sky130_fd_sc_hd__and3_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _09673_/X _09675_/X _09778_/C _09767_/A VGND VGND VPWR VPWR _09679_/C sky130_fd_sc_hd__a2bb2o_1
X_06889_ _07962_/B VGND VGND VPWR VPWR _07968_/B sky130_fd_sc_hd__buf_2
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ _13447_/Q _09450_/B VGND VGND VPWR VPWR _08630_/A sky130_fd_sc_hd__xnor2_1
XFILLER_27_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _13441_/Q _09417_/B VGND VGND VPWR VPWR _08572_/A sky130_fd_sc_hd__and2_1
XFILLER_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11570_ _13643_/Q _11574_/B VGND VGND VPWR VPWR _11571_/A sky130_fd_sc_hd__and2_1
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10521_ _10555_/B _10521_/B VGND VGND VPWR VPWR _10533_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13240_ _14010_/CLK _13240_/D VGND VGND VPWR VPWR _13512_/D sky130_fd_sc_hd__dfxtp_1
X_10452_ _10452_/A _10452_/B VGND VGND VPWR VPWR _10453_/B sky130_fd_sc_hd__xnor2_1
XFILLER_10_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13171_ _13666_/CLK _13171_/D VGND VGND VPWR VPWR _13171_/Q sky130_fd_sc_hd__dfxtp_2
X_10383_ _13517_/Q _13518_/Q _10387_/B _10382_/X VGND VGND VPWR VPWR _10393_/A sky130_fd_sc_hd__a31o_1
XFILLER_151_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12122_ _14476_/Q _11988_/X _12128_/S VGND VGND VPWR VPWR _12123_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12053_ _12053_/A VGND VGND VPWR VPWR _14445_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11004_ _10932_/X _11001_/Y _11003_/Y _10946_/X VGND VGND VPWR VPWR _11005_/B sky130_fd_sc_hd__a211o_1
Xclkbuf_3_6_0_clk clkbuf_3_7_0_clk/A VGND VGND VPWR VPWR clkbuf_3_6_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12955_ _13039_/CLK hold252/X VGND VGND VPWR VPWR _12955_/Q sky130_fd_sc_hd__dfxtp_1
X_11906_ _11906_/A VGND VGND VPWR VPWR _14260_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12886_ _12930_/CLK _12886_/D hold1/X VGND VGND VPWR VPWR _12886_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ _11837_/A VGND VGND VPWR VPWR _14166_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14625_ _14633_/CLK _14625_/D VGND VGND VPWR VPWR _14625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _14557_/CLK _14556_/D VGND VGND VPWR VPWR _14556_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _13557_/Q _11772_/B VGND VGND VPWR VPWR _11769_/A sky130_fd_sc_hd__and2_1
XFILLER_119_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13507_ _13811_/CLK hold18/X VGND VGND VPWR VPWR _13507_/Q sky130_fd_sc_hd__dfxtp_1
X_10719_ _10719_/A VGND VGND VPWR VPWR _12937_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14487_ _14619_/CLK _14487_/D VGND VGND VPWR VPWR _14487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11699_ _11699_/A VGND VGND VPWR VPWR _14031_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13438_ _13476_/CLK _13438_/D repeater56/X VGND VGND VPWR VPWR _13438_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_127_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13369_ _13621_/CLK _13369_/D repeater56/X VGND VGND VPWR VPWR _13369_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07930_ _07939_/A _07930_/B VGND VGND VPWR VPWR _07949_/B sky130_fd_sc_hd__nand2_1
XFILLER_111_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07861_ _06781_/B _07860_/X _07861_/S VGND VGND VPWR VPWR _07862_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09600_ _09600_/A VGND VGND VPWR VPWR _09609_/S sky130_fd_sc_hd__clkbuf_2
X_06812_ _06863_/A _06812_/B VGND VGND VPWR VPWR _06813_/C sky130_fd_sc_hd__nor2_2
X_07792_ _07780_/Y _07791_/Y _07800_/S VGND VGND VPWR VPWR _07793_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09531_ _09532_/A _09532_/B _09532_/C VGND VGND VPWR VPWR _09531_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06743_ _06743_/A _06743_/B VGND VGND VPWR VPWR _06743_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09462_ _08504_/X _09461_/Y _08642_/X VGND VGND VPWR VPWR _13602_/D sky130_fd_sc_hd__a21o_1
X_06674_ _06746_/S _13342_/Q _06674_/C VGND VGND VPWR VPWR _06674_/X sky130_fd_sc_hd__and3b_1
XFILLER_36_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08413_ _08413_/A VGND VGND VPWR VPWR _12737_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09393_ _08784_/X _09419_/A _09392_/X _08515_/X VGND VGND VPWR VPWR _13593_/D sky130_fd_sc_hd__a31o_1
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08344_ _13385_/Q _08340_/X _08157_/X VGND VGND VPWR VPWR _08344_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08275_ _08256_/A _08257_/A _08256_/B _08267_/A _08274_/X VGND VGND VPWR VPWR _08276_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_164_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07226_ _13170_/Q VGND VGND VPWR VPWR _07299_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_118_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07157_ _07136_/Y _07156_/Y _07199_/S VGND VGND VPWR VPWR _07158_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06108_ _06108_/A VGND VGND VPWR VPWR _13944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07088_ _07106_/A _07106_/B VGND VGND VPWR VPWR _07107_/A sky130_fd_sc_hd__xnor2_1
XFILLER_160_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06039_ input17/X hold42/A _06035_/A VGND VGND VPWR VPWR _06041_/A sky130_fd_sc_hd__o21a_1
XFILLER_154_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09729_ _09722_/B _09726_/X _09774_/S VGND VGND VPWR VPWR _09730_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12740_ _14696_/CLK _12740_/D VGND VGND VPWR VPWR hold109/A sky130_fd_sc_hd__dfxtp_1
XFILLER_83_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12671_ _14439_/CLK _12671_/D VGND VGND VPWR VPWR _12671_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14410_/CLK _14410_/D VGND VGND VPWR VPWR hold94/A sky130_fd_sc_hd__dfxtp_2
X_11622_ _11622_/A VGND VGND VPWR VPWR _13987_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14341_ _14697_/CLK hold484/X VGND VGND VPWR VPWR _14341_/Q sky130_fd_sc_hd__dfxtp_1
X_11553_ _11553_/A VGND VGND VPWR VPWR _13859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10504_ _10438_/B _10439_/A _10441_/A VGND VGND VPWR VPWR _10504_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_11_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14272_ _14720_/CLK _14272_/D VGND VGND VPWR VPWR _14272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11484_ _11484_/A VGND VGND VPWR VPWR _13829_/D sky130_fd_sc_hd__clkbuf_1
X_13223_ _13606_/CLK hold147/X VGND VGND VPWR VPWR _13223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10435_ _10444_/B VGND VGND VPWR VPWR _10439_/A sky130_fd_sc_hd__inv_2
XFILLER_136_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13154_ _13377_/CLK _13154_/D repeater57/X VGND VGND VPWR VPWR _13154_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10366_ _10432_/A _10366_/B _10378_/A VGND VGND VPWR VPWR _10367_/A sky130_fd_sc_hd__and3_1
XFILLER_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _12105_/A VGND VGND VPWR VPWR _14468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13085_ _13565_/CLK hold365/X VGND VGND VPWR VPWR _13085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10297_ hold118/X hold41/X _10296_/X VGND VGND VPWR VPWR _13814_/D sky130_fd_sc_hd__o21a_1
X_12036_ _12678_/Q _12036_/B VGND VGND VPWR VPWR _12037_/A sky130_fd_sc_hd__and2_1
XFILLER_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13987_ _14357_/CLK _13987_/D VGND VGND VPWR VPWR _13987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _12970_/CLK _12938_/D VGND VGND VPWR VPWR hold143/A sky130_fd_sc_hd__dfxtp_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _13811_/CLK _12869_/D VGND VGND VPWR VPWR hold323/A sky130_fd_sc_hd__dfxtp_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14608_ _14608_/CLK _14608_/D VGND VGND VPWR VPWR _14608_/Q sky130_fd_sc_hd__dfxtp_1
X_06390_ _10679_/A _06622_/B VGND VGND VPWR VPWR _06391_/B sky130_fd_sc_hd__nand2_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14539_ _14539_/CLK _14539_/D VGND VGND VPWR VPWR _14539_/Q sky130_fd_sc_hd__dfxtp_1
X_08060_ _12967_/Q _13267_/Q _08062_/S VGND VGND VPWR VPWR _08061_/A sky130_fd_sc_hd__mux2_1
X_07011_ _14634_/Q VGND VGND VPWR VPWR _07031_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08962_ _08962_/A _08962_/B VGND VGND VPWR VPWR _08966_/B sky130_fd_sc_hd__and2_1
X_07913_ _07914_/A _07914_/B _07916_/B VGND VGND VPWR VPWR _07913_/X sky130_fd_sc_hd__a21o_1
X_08893_ _08893_/A VGND VGND VPWR VPWR _14249_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07844_ _07844_/A VGND VGND VPWR VPWR _13258_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07775_ _07787_/A _07787_/B _07760_/A VGND VGND VPWR VPWR _07776_/B sky130_fd_sc_hd__a21oi_1
XFILLER_83_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09514_ _09508_/Y _09510_/X _09534_/A VGND VGND VPWR VPWR _09514_/X sky130_fd_sc_hd__a21o_1
XFILLER_25_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06726_ _13003_/Q _07840_/B VGND VGND VPWR VPWR _06727_/B sky130_fd_sc_hd__nor2_1
XFILLER_65_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09445_ _09443_/A _09448_/C _09448_/D VGND VGND VPWR VPWR _09455_/B sky130_fd_sc_hd__o21ba_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06657_ _12999_/Q _06690_/A _07804_/C VGND VGND VPWR VPWR _06659_/A sky130_fd_sc_hd__and3_1
XFILLER_52_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09376_ _13591_/Q _09383_/B VGND VGND VPWR VPWR _09377_/C sky130_fd_sc_hd__nand2_1
X_06588_ _12896_/Q _06595_/B VGND VGND VPWR VPWR _06590_/A sky130_fd_sc_hd__and2_1
XFILLER_149_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08327_ _13378_/Q _13379_/Q _08325_/D _13380_/Q VGND VGND VPWR VPWR _08328_/C sky130_fd_sc_hd__a31o_1
XFILLER_149_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08258_ _08252_/B _08257_/Y _08286_/S VGND VGND VPWR VPWR _08259_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07209_ _07209_/A _07209_/B VGND VGND VPWR VPWR _07209_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_4_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08189_ _08189_/A _08189_/B VGND VGND VPWR VPWR _08193_/A sky130_fd_sc_hd__or2_1
X_10220_ _14099_/Q _14083_/Q _10224_/S VGND VGND VPWR VPWR _10221_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10151_ _14285_/D _10150_/X _14294_/D VGND VGND VPWR VPWR _10151_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10082_ _10073_/X _10081_/X _14049_/D VGND VGND VPWR VPWR _10082_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13910_ _13978_/CLK _13910_/D VGND VGND VPWR VPWR _13910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13841_ _14725_/CLK _13841_/D VGND VGND VPWR VPWR _13841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13772_ _14275_/CLK _13772_/D VGND VGND VPWR VPWR _13772_/Q sky130_fd_sc_hd__dfxtp_1
X_10984_ _14599_/Q _14561_/Q _14492_/Q _14444_/Q _10969_/X _10970_/X VGND VGND VPWR
+ VPWR _10985_/A sky130_fd_sc_hd__mux4_1
X_12723_ _13606_/CLK _12723_/D VGND VGND VPWR VPWR hold465/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12654_ _14082_/CLK hold496/X _12609_/A VGND VGND VPWR VPWR hold501/A sky130_fd_sc_hd__dfrtp_1
XFILLER_90_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11605_ _11605_/A VGND VGND VPWR VPWR _13979_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12585_ _12585_/A _14730_/Q VGND VGND VPWR VPWR _12585_/X sky130_fd_sc_hd__or2_1
XFILLER_157_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14324_ _14688_/CLK _14324_/D VGND VGND VPWR VPWR _14324_/Q sky130_fd_sc_hd__dfxtp_1
X_11536_ _11536_/A VGND VGND VPWR VPWR _13851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14255_ _14256_/CLK _14255_/D VGND VGND VPWR VPWR _14255_/Q sky130_fd_sc_hd__dfxtp_1
X_11467_ _13824_/Q _11465_/X _11479_/S VGND VGND VPWR VPWR _11468_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13206_ _14012_/CLK hold224/X VGND VGND VPWR VPWR _13206_/Q sky130_fd_sc_hd__dfxtp_1
X_10418_ _10417_/B _10418_/B VGND VGND VPWR VPWR _10419_/B sky130_fd_sc_hd__and2b_1
X_14186_ _14201_/CLK _14186_/D VGND VGND VPWR VPWR _14186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11398_ _11398_/A VGND VGND VPWR VPWR _13791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13137_ _13359_/CLK _13137_/D hold1/X VGND VGND VPWR VPWR _13137_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10349_ _10349_/A _13121_/D VGND VGND VPWR VPWR _10352_/A sky130_fd_sc_hd__xnor2_1
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _14555_/CLK _13068_/D VGND VGND VPWR VPWR hold446/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12019_ _12019_/A VGND VGND VPWR VPWR _12019_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07560_ _09258_/B VGND VGND VPWR VPWR _09250_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_81_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06511_ _06513_/B _06554_/C VGND VGND VPWR VPWR _06514_/B sky130_fd_sc_hd__and2_1
X_07491_ _07498_/A _07491_/B VGND VGND VPWR VPWR _07504_/C sky130_fd_sc_hd__nand2_1
XFILLER_34_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09230_ _09230_/A _09242_/C VGND VGND VPWR VPWR _09230_/Y sky130_fd_sc_hd__xnor2_1
X_06442_ _14435_/Q _14433_/Q _06458_/S VGND VGND VPWR VPWR _06442_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09161_ _09161_/A _09161_/B _09161_/C VGND VGND VPWR VPWR _09161_/X sky130_fd_sc_hd__or3_1
X_06373_ _13389_/D hold41/A _13388_/D VGND VGND VPWR VPWR _06373_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08112_ _08296_/B _13354_/Q VGND VGND VPWR VPWR _08113_/B sky130_fd_sc_hd__nand2_1
X_09092_ _09089_/B _09089_/C _09089_/A VGND VGND VPWR VPWR _09095_/A sky130_fd_sc_hd__o21ba_1
X_08043_ _12959_/Q _13259_/Q _08051_/S VGND VGND VPWR VPWR _08044_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09994_ _10636_/A _14626_/Q VGND VGND VPWR VPWR _09994_/X sky130_fd_sc_hd__and2b_1
X_08945_ _08924_/Y _08944_/Y _08987_/S VGND VGND VPWR VPWR _08946_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08876_ _08894_/A _08894_/B VGND VGND VPWR VPWR _08895_/A sky130_fd_sc_hd__xnor2_1
XFILLER_151_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07827_ _13255_/Q _07819_/B _07815_/A _07815_/B _07821_/X VGND VGND VPWR VPWR _07828_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_57_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07758_ _07732_/A _07732_/B _07757_/X VGND VGND VPWR VPWR _07759_/C sky130_fd_sc_hd__a21oi_1
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06709_ _06710_/B VGND VGND VPWR VPWR _07832_/B sky130_fd_sc_hd__clkbuf_2
X_07689_ _07689_/A _07689_/B _07689_/C VGND VGND VPWR VPWR _07705_/B sky130_fd_sc_hd__or3_1
XFILLER_44_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09428_ _09447_/C _09454_/A _09427_/X VGND VGND VPWR VPWR _09428_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_157_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09359_ _13315_/Q _13553_/Q _10822_/A VGND VGND VPWR VPWR _09360_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12370_ _12370_/A VGND VGND VPWR VPWR _14607_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11321_ _13767_/Q _11320_/X _11327_/S VGND VGND VPWR VPWR _11322_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14040_ _14042_/CLK _14040_/D VGND VGND VPWR VPWR _14040_/Q sky130_fd_sc_hd__dfxtp_1
X_11252_ _10944_/A _11249_/Y _11251_/Y _10929_/A VGND VGND VPWR VPWR _11253_/B sky130_fd_sc_hd__a211o_1
XFILLER_134_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10203_ _14402_/Q _14394_/Q _10627_/A VGND VGND VPWR VPWR _10203_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11183_ _11183_/A _11155_/X VGND VGND VPWR VPWR _11183_/X sky130_fd_sc_hd__or2b_1
XFILLER_122_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10134_ _10134_/A VGND VGND VPWR VPWR _14181_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10065_ _14043_/D _10064_/X _10092_/S VGND VGND VPWR VPWR _10066_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13824_ _14536_/CLK _13824_/D VGND VGND VPWR VPWR _13824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10967_ _12645_/A _10964_/X _10966_/X _10929_/X VGND VGND VPWR VPWR _10967_/X sky130_fd_sc_hd__o211a_1
X_13755_ _14703_/CLK _13755_/D VGND VGND VPWR VPWR _13755_/Q sky130_fd_sc_hd__dfxtp_1
X_12706_ _14108_/CLK _12706_/D VGND VGND VPWR VPWR hold290/A sky130_fd_sc_hd__dfxtp_1
X_10898_ _14747_/Q _14737_/Q VGND VGND VPWR VPWR _10899_/D sky130_fd_sc_hd__xor2_1
X_13686_ _13686_/CLK _13686_/D repeater56/X VGND VGND VPWR VPWR _13686_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12637_ _12637_/A _12637_/B VGND VGND VPWR VPWR _14743_/D sky130_fd_sc_hd__nor2_1
XFILLER_31_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12568_ _14744_/Q VGND VGND VPWR VPWR _12568_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14307_ _14602_/CLK _14307_/D VGND VGND VPWR VPWR _14307_/Q sky130_fd_sc_hd__dfxtp_1
X_11519_ _12022_/A VGND VGND VPWR VPWR _11519_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12499_ _12499_/A VGND VGND VPWR VPWR _14679_/D sky130_fd_sc_hd__clkbuf_1
Xhold207 hold207/A VGND VGND VPWR VPWR hold207/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold218 hold218/A VGND VGND VPWR VPWR hold218/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold229 hold229/A VGND VGND VPWR VPWR hold229/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14238_ _14510_/CLK _14238_/D VGND VGND VPWR VPWR _14238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14169_ _14196_/CLK _14169_/D VGND VGND VPWR VPWR _14169_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ _13027_/Q _08008_/B VGND VGND VPWR VPWR _06991_/X sky130_fd_sc_hd__or2_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08730_ _13457_/Q _08730_/B VGND VGND VPWR VPWR _08731_/B sky130_fd_sc_hd__nor2_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05942_ _13871_/Q _13872_/Q _13873_/Q _13874_/Q VGND VGND VPWR VPWR _05944_/B sky130_fd_sc_hd__or4_1
XFILLER_38_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08661_ _13450_/Q _09472_/B VGND VGND VPWR VPWR _08662_/B sky130_fd_sc_hd__nor2_1
XFILLER_82_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07612_ _07668_/C VGND VGND VPWR VPWR _07723_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08592_ _09424_/B _09424_/C VGND VGND VPWR VPWR _08592_/X sky130_fd_sc_hd__and2_1
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07543_ _07547_/B _07543_/B VGND VGND VPWR VPWR _07543_/X sky130_fd_sc_hd__xor2_1
X_07474_ _09215_/A VGND VGND VPWR VPWR _07499_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09213_ _09214_/A _09214_/B _09220_/D VGND VGND VPWR VPWR _09213_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06425_ _14438_/Q _14436_/Q _06425_/S VGND VGND VPWR VPWR _06425_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09144_ _08157_/X _09140_/B _09142_/Y _09143_/X VGND VGND VPWR VPWR _13532_/D sky130_fd_sc_hd__a22o_1
X_06356_ _06355_/Y _06025_/B _14590_/D _14682_/Q VGND VGND VPWR VPWR _12875_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_136_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09075_ _13235_/Q _13464_/Q _09075_/S VGND VGND VPWR VPWR _09076_/A sky130_fd_sc_hd__mux2_1
X_06287_ hold52/A _13952_/D _06287_/C _06287_/D VGND VGND VPWR VPWR hold503/A sky130_fd_sc_hd__nand4_1
XFILLER_107_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08026_ _12952_/Q _13252_/Q _10818_/B VGND VGND VPWR VPWR _08027_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09977_ _10597_/A _14592_/Q VGND VGND VPWR VPWR _09977_/X sky130_fd_sc_hd__and2b_1
XFILLER_89_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08928_ _08951_/A _08978_/A _08951_/B _08929_/A VGND VGND VPWR VPWR _08930_/A sky130_fd_sc_hd__a22oi_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08859_ _08860_/A _08860_/B VGND VGND VPWR VPWR _08861_/A sky130_fd_sc_hd__and2_1
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _11870_/A VGND VGND VPWR VPWR _14232_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ _10821_/A VGND VGND VPWR VPWR _13072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13540_ _13558_/CLK _13540_/D _12609_/A VGND VGND VPWR VPWR _13540_/Q sky130_fd_sc_hd__dfrtp_2
X_10752_ _10752_/A VGND VGND VPWR VPWR _13040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13471_ _13476_/CLK _13471_/D VGND VGND VPWR VPWR _13471_/Q sky130_fd_sc_hd__dfxtp_1
X_10683_ _12878_/Q _10687_/B VGND VGND VPWR VPWR _10684_/A sky130_fd_sc_hd__and2_1
X_12422_ _12484_/A _12484_/B input5/X VGND VGND VPWR VPWR _12423_/A sky130_fd_sc_hd__and3_1
XFILLER_40_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12353_ _14600_/Q _11965_/X _12353_/S VGND VGND VPWR VPWR _12354_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11304_ _14701_/Q VGND VGND VPWR VPWR _11304_/X sky130_fd_sc_hd__buf_2
XFILLER_154_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12284_ _12284_/A VGND VGND VPWR VPWR _14558_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14023_ _14713_/CLK _14023_/D VGND VGND VPWR VPWR _14023_/Q sky130_fd_sc_hd__dfxtp_1
X_11235_ _11235_/A _10960_/A VGND VGND VPWR VPWR _11235_/X sky130_fd_sc_hd__or2b_1
XFILLER_122_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11166_ _11166_/A VGND VGND VPWR VPWR _11166_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10117_ _10616_/D _10116_/X _10119_/S VGND VGND VPWR VPWR _10118_/A sky130_fd_sc_hd__mux2_1
X_11097_ _11108_/A _11097_/B VGND VGND VPWR VPWR _11097_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10048_ _13804_/Q _13788_/Q _10050_/S VGND VGND VPWR VPWR _10049_/A sky130_fd_sc_hd__mux2_1
Xhold90 hold90/A VGND VGND VPWR VPWR hold90/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_152_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13807_ _13811_/CLK _13807_/D VGND VGND VPWR VPWR _13807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11999_ _11999_/A VGND VGND VPWR VPWR _14309_/D sky130_fd_sc_hd__clkbuf_1
X_13738_ _13963_/CLK hold172/X VGND VGND VPWR VPWR _13738_/Q sky130_fd_sc_hd__dfxtp_1
X_13669_ _14251_/CLK _13669_/D repeater56/X VGND VGND VPWR VPWR _13669_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06210_ _14405_/Q _14397_/Q hold94/A VGND VGND VPWR VPWR _06215_/C sky130_fd_sc_hd__mux2_1
X_07190_ _07190_/A _07190_/B _07203_/C _07190_/D VGND VGND VPWR VPWR _07191_/B sky130_fd_sc_hd__and4_1
XFILLER_129_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06141_ _14189_/Q _14181_/Q _14194_/D VGND VGND VPWR VPWR _06145_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06072_ _13962_/D VGND VGND VPWR VPWR _06256_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_144_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09900_ _13697_/Q _09886_/A _09893_/B _13698_/Q VGND VGND VPWR VPWR _09901_/B sky130_fd_sc_hd__a31o_1
XFILLER_104_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09831_ _09812_/A _09822_/A _09822_/B VGND VGND VPWR VPWR _09831_/X sky130_fd_sc_hd__o21ba_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06974_ _07940_/A VGND VGND VPWR VPWR _06974_/X sky130_fd_sc_hd__buf_2
XFILLER_86_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09762_ _09753_/A _09753_/B _09749_/A VGND VGND VPWR VPWR _09763_/B sky130_fd_sc_hd__o21bai_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05925_ _13740_/Q _13741_/Q _13742_/Q _13743_/Q VGND VGND VPWR VPWR _05928_/A sky130_fd_sc_hd__and4_1
X_08713_ _08713_/A _08713_/B VGND VGND VPWR VPWR _08741_/A sky130_fd_sc_hd__nand2_1
X_09693_ _09682_/A _09680_/X _09681_/A VGND VGND VPWR VPWR _09697_/A sky130_fd_sc_hd__a21o_1
XFILLER_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08644_ _08644_/A _08644_/B VGND VGND VPWR VPWR _08654_/A sky130_fd_sc_hd__nor2_1
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _08622_/A _08574_/B _08542_/A VGND VGND VPWR VPWR _08575_/Y sky130_fd_sc_hd__a21oi_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07526_ _09215_/A VGND VGND VPWR VPWR _07526_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07457_ _13143_/Q _09163_/B _07438_/A VGND VGND VPWR VPWR _07457_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06408_ _10679_/A _06391_/A _06399_/B _06397_/X VGND VGND VPWR VPWR _06421_/A sky130_fd_sc_hd__a31o_1
XFILLER_10_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07388_ _07400_/A _07388_/B VGND VGND VPWR VPWR _07389_/B sky130_fd_sc_hd__nor2_1
X_09127_ _13529_/Q _07356_/B _09122_/X VGND VGND VPWR VPWR _09128_/B sky130_fd_sc_hd__a21bo_1
X_06339_ _14106_/Q _14090_/Q _06341_/S VGND VGND VPWR VPWR _06340_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09058_ _13227_/Q _13456_/Q _09064_/S VGND VGND VPWR VPWR _09059_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08009_ _08003_/A _08004_/Y _08007_/Y _08008_/X VGND VGND VPWR VPWR _08009_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_135_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11020_ _11162_/A VGND VGND VPWR VPWR _11020_/X sky130_fd_sc_hd__buf_2
XFILLER_106_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12971_ _13273_/CLK hold143/X VGND VGND VPWR VPWR _12971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14710_ _14710_/CLK _14710_/D VGND VGND VPWR VPWR _14710_/Q sky130_fd_sc_hd__dfxtp_1
X_11922_ _11922_/A VGND VGND VPWR VPWR _14267_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _14643_/CLK _14641_/D VGND VGND VPWR VPWR _14641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _14225_/Q _11462_/X _11853_/S VGND VGND VPWR VPWR _11854_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _13022_/Q _10812_/B VGND VGND VPWR VPWR _10805_/A sky130_fd_sc_hd__and2_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14572_ _14610_/CLK _14572_/D VGND VGND VPWR VPWR _14572_/Q sky130_fd_sc_hd__dfxtp_1
X_11784_ _13564_/Q _11784_/B VGND VGND VPWR VPWR _11785_/A sky130_fd_sc_hd__and2_1
XFILLER_158_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13523_ _13525_/CLK _13523_/D hold1/X VGND VGND VPWR VPWR _13523_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_40_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10735_ _10735_/A VGND VGND VPWR VPWR _12944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10666_ _14339_/Q _14340_/Q _10666_/C VGND VGND VPWR VPWR _10671_/C sky130_fd_sc_hd__and3_1
X_13454_ _13605_/CLK _13454_/D repeater57/X VGND VGND VPWR VPWR _13454_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12405_ _12405_/A VGND VGND VPWR VPWR _14634_/D sky130_fd_sc_hd__clkbuf_1
X_13385_ _14530_/CLK _13385_/D _12609_/A VGND VGND VPWR VPWR _13385_/Q sky130_fd_sc_hd__dfrtp_1
X_10597_ _10597_/A _14629_/Q VGND VGND VPWR VPWR _14622_/D sky130_fd_sc_hd__xor2_1
XFILLER_154_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12336_ _14640_/Q _12340_/B _12336_/C VGND VGND VPWR VPWR _12337_/A sky130_fd_sc_hd__and3_1
XFILLER_99_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12267_ _12267_/A VGND VGND VPWR VPWR _14548_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11218_ _11159_/X _11215_/Y _11217_/Y _11166_/X VGND VGND VPWR VPWR _11219_/B sky130_fd_sc_hd__a211o_1
X_14006_ _14679_/CLK _14006_/D VGND VGND VPWR VPWR _14006_/Q sky130_fd_sc_hd__dfxtp_1
X_12198_ _14510_/Q _12019_/X _12202_/S VGND VGND VPWR VPWR _12199_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11149_ _13332_/Q _11079_/X _11142_/X _11148_/Y VGND VGND VPWR VPWR _13332_/D sky130_fd_sc_hd__o22a_1
XFILLER_95_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06690_ _06690_/A _06690_/B _06689_/X VGND VGND VPWR VPWR _06786_/A sky130_fd_sc_hd__nor3b_2
XFILLER_24_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08360_ _13078_/Q _13359_/Q _08362_/S VGND VGND VPWR VPWR _08361_/A sky130_fd_sc_hd__mux2_1
X_07311_ _07311_/A _07311_/B _07311_/C VGND VGND VPWR VPWR _07349_/A sky130_fd_sc_hd__and3_1
X_08291_ _13370_/Q _08294_/A _08157_/X VGND VGND VPWR VPWR _08291_/Y sky130_fd_sc_hd__a21oi_1
X_07242_ _13666_/Q _13664_/Q _13170_/Q VGND VGND VPWR VPWR _07428_/B sky130_fd_sc_hd__mux2_1
XFILLER_158_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07173_ _07174_/A _07174_/B VGND VGND VPWR VPWR _07178_/A sky130_fd_sc_hd__nor2_1
XFILLER_118_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06124_ _06124_/A VGND VGND VPWR VPWR _14149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14753__64 VGND VGND VPWR VPWR _14753__64/HI data_o[27] sky130_fd_sc_hd__conb_1
XFILLER_132_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06055_ _13977_/Q VGND VGND VPWR VPWR _10020_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_160_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09814_ _09795_/A _09804_/Y _09795_/B _09803_/A _09792_/A VGND VGND VPWR VPWR _09815_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_143_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09745_ _09735_/A _14220_/Q _09836_/B _09778_/A VGND VGND VPWR VPWR _09746_/C sky130_fd_sc_hd__a31o_1
X_06957_ _06968_/A _06967_/A _06976_/A VGND VGND VPWR VPWR _06957_/X sky130_fd_sc_hd__o21a_1
XFILLER_27_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05908_ _13803_/Q _13804_/Q _13805_/Q _13806_/Q VGND VGND VPWR VPWR _05909_/C sky130_fd_sc_hd__and4_1
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06888_ _06899_/A _06924_/A VGND VGND VPWR VPWR _06888_/Y sky130_fd_sc_hd__xnor2_1
X_09676_ _14440_/Q _14219_/Q _14217_/Q _14215_/Q _09688_/S _13710_/Q VGND VGND VPWR
+ VPWR _09778_/C sky130_fd_sc_hd__mux4_2
XFILLER_54_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _09451_/B VGND VGND VPWR VPWR _09450_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08558_ _08558_/A _08572_/B VGND VGND VPWR VPWR _08561_/A sky130_fd_sc_hd__or2_1
XFILLER_11_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07509_ _07532_/A _07510_/B VGND VGND VPWR VPWR _07509_/X sky130_fd_sc_hd__or2_1
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08489_ _08434_/Y _08606_/B _08488_/X _08431_/X VGND VGND VPWR VPWR _08489_/X sky130_fd_sc_hd__a22o_1
XFILLER_11_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10520_ _10520_/A _10539_/A VGND VGND VPWR VPWR _10525_/A sky130_fd_sc_hd__or2_1
XFILLER_10_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10451_ hold186/A _10449_/A _10444_/B VGND VGND VPWR VPWR _10452_/B sky130_fd_sc_hd__o21ai_1
XFILLER_109_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13170_ _13666_/CLK _13170_/D VGND VGND VPWR VPWR _13170_/Q sky130_fd_sc_hd__dfxtp_1
X_10382_ _14211_/D _13516_/Q _13519_/Q _13520_/Q VGND VGND VPWR VPWR _10382_/X sky130_fd_sc_hd__and4_1
XFILLER_164_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12121_ _12121_/A VGND VGND VPWR VPWR _14475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12052_ _11294_/X _14445_/Q _12052_/S VGND VGND VPWR VPWR _12053_/A sky130_fd_sc_hd__mux2_1
Xhold390 hold390/A VGND VGND VPWR VPWR hold390/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11003_ _11035_/A _11003_/B VGND VGND VPWR VPWR _11003_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12954_ _13039_/CLK hold234/X VGND VGND VPWR VPWR _12954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11905_ _14260_/Q _11459_/X _11907_/S VGND VGND VPWR VPWR _11906_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _12885_/CLK _12885_/D hold1/X VGND VGND VPWR VPWR _12885_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _14636_/CLK _14629_/Q VGND VGND VPWR VPWR _14624_/Q sky130_fd_sc_hd__dfxtp_1
X_11836_ _12679_/Q _11836_/B VGND VGND VPWR VPWR _11837_/A sky130_fd_sc_hd__and2_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14555_ _14555_/CLK _14555_/D VGND VGND VPWR VPWR hold120/A sky130_fd_sc_hd__dfxtp_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _11767_/A VGND VGND VPWR VPWR _14074_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13506_ _13698_/CLK hold397/X VGND VGND VPWR VPWR hold456/A sky130_fd_sc_hd__dfxtp_1
X_10718_ _12894_/Q _10720_/B VGND VGND VPWR VPWR _10719_/A sky130_fd_sc_hd__and2_1
X_14486_ _14617_/CLK _14486_/D VGND VGND VPWR VPWR _14486_/Q sky130_fd_sc_hd__dfxtp_1
X_11698_ _14031_/Q _11507_/X _11700_/S VGND VGND VPWR VPWR _11699_/A sky130_fd_sc_hd__mux2_1
X_13437_ _13593_/CLK _13437_/D repeater56/X VGND VGND VPWR VPWR _13437_/Q sky130_fd_sc_hd__dfrtp_1
X_10649_ _13556_/Q _11772_/B VGND VGND VPWR VPWR _10650_/A sky130_fd_sc_hd__and2_1
X_13368_ _13423_/CLK _13368_/D repeater57/X VGND VGND VPWR VPWR _13368_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12319_ _12319_/A VGND VGND VPWR VPWR _14574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13299_ _13303_/CLK hold459/X VGND VGND VPWR VPWR _13299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07860_ _07860_/A _07860_/B VGND VGND VPWR VPWR _07860_/X sky130_fd_sc_hd__xor2_1
XFILLER_96_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06811_ _06811_/A VGND VGND VPWR VPWR _06813_/B sky130_fd_sc_hd__inv_2
X_07791_ _07791_/A _07791_/B VGND VGND VPWR VPWR _07791_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_95_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09530_ _13612_/Q _09530_/B VGND VGND VPWR VPWR _09532_/C sky130_fd_sc_hd__xor2_1
X_06742_ _06727_/B _06731_/B _06739_/Y _06725_/A VGND VGND VPWR VPWR _06743_/B sky130_fd_sc_hd__o211a_1
XFILLER_36_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09461_ _09478_/A _09466_/B VGND VGND VPWR VPWR _09461_/Y sky130_fd_sc_hd__xnor2_1
X_06673_ _13037_/Q VGND VGND VPWR VPWR _06746_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_184_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _14749_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08412_ hold469/X _13382_/Q _08418_/S VGND VGND VPWR VPWR _08413_/A sky130_fd_sc_hd__mux2_1
X_09392_ _09382_/A _09390_/X _09391_/B VGND VGND VPWR VPWR _09392_/X sky130_fd_sc_hd__a21bo_1
XFILLER_33_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08343_ _08343_/A VGND VGND VPWR VPWR _13384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08274_ _08253_/A _08265_/A _08265_/B VGND VGND VPWR VPWR _08274_/X sky130_fd_sc_hd__o21ba_1
XFILLER_138_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07225_ _13171_/Q VGND VGND VPWR VPWR _07266_/A sky130_fd_sc_hd__inv_2
XFILLER_164_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07156_ _07156_/A _07156_/B VGND VGND VPWR VPWR _07156_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06107_ _13798_/Q _12680_/Q _10050_/S VGND VGND VPWR VPWR _06108_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07087_ _07087_/A _07114_/B VGND VGND VPWR VPWR _07106_/B sky130_fd_sc_hd__nor2_1
XFILLER_160_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06038_ hold41/A VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__inv_2
XFILLER_59_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07989_ _13278_/Q _07989_/B VGND VGND VPWR VPWR _07990_/B sky130_fd_sc_hd__or2_1
XFILLER_68_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09728_ _09855_/A VGND VGND VPWR VPWR _09774_/S sky130_fd_sc_hd__buf_2
XFILLER_90_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_175_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _14600_/CLK sky130_fd_sc_hd__clkbuf_16
X_09659_ _09758_/A VGND VGND VPWR VPWR _09778_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12670_ _13351_/CLK _12670_/D VGND VGND VPWR VPWR _12992_/D sky130_fd_sc_hd__dfxtp_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11621_ _13987_/Q _11475_/X _11623_/S VGND VGND VPWR VPWR _11622_/A sky130_fd_sc_hd__mux2_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14340_ _14697_/CLK hold491/X VGND VGND VPWR VPWR _14340_/Q sky130_fd_sc_hd__dfxtp_1
X_11552_ _13635_/Q _11552_/B VGND VGND VPWR VPWR _11553_/A sky130_fd_sc_hd__and2_1
XFILLER_11_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10503_ _10503_/A _10503_/B VGND VGND VPWR VPWR _13477_/D sky130_fd_sc_hd__nand2_1
XFILLER_156_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14271_ _14716_/CLK _14271_/D VGND VGND VPWR VPWR _14271_/Q sky130_fd_sc_hd__dfxtp_1
X_11483_ _13829_/Q _11481_/X _11495_/S VGND VGND VPWR VPWR _11484_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10434_ _10485_/A VGND VGND VPWR VPWR _10444_/B sky130_fd_sc_hd__clkbuf_2
X_13222_ _13606_/CLK hold405/X VGND VGND VPWR VPWR _13222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10365_ _10386_/A _10376_/A VGND VGND VPWR VPWR _10378_/A sky130_fd_sc_hd__nand2_1
X_13153_ _13552_/CLK _13153_/D _12609_/A VGND VGND VPWR VPWR _13153_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _14468_/Q _11962_/X _12106_/S VGND VGND VPWR VPWR _12105_/A sky130_fd_sc_hd__mux2_1
X_13084_ _13528_/CLK hold126/X VGND VGND VPWR VPWR _13084_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10296_ hold42/X _10296_/B VGND VGND VPWR VPWR _10296_/X sky130_fd_sc_hd__or2_1
XFILLER_3_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12035_ _12035_/A VGND VGND VPWR VPWR _14326_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13986_ _14710_/CLK _13986_/D VGND VGND VPWR VPWR _13986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12937_ _12970_/CLK _12937_/D VGND VGND VPWR VPWR hold321/A sky130_fd_sc_hd__dfxtp_1
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_166_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _14357_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _13811_/CLK _12868_/D VGND VGND VPWR VPWR hold388/A sky130_fd_sc_hd__dfxtp_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14607_ _14717_/CLK _14607_/D VGND VGND VPWR VPWR _14607_/Q sky130_fd_sc_hd__dfxtp_1
X_11819_ _11819_/A VGND VGND VPWR VPWR _11828_/B sky130_fd_sc_hd__clkbuf_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _14275_/CLK _12799_/D VGND VGND VPWR VPWR hold349/A sky130_fd_sc_hd__dfxtp_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14538_ _14697_/CLK _14538_/D VGND VGND VPWR VPWR _14538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14469_ _14705_/CLK _14469_/D VGND VGND VPWR VPWR _14469_/Q sky130_fd_sc_hd__dfxtp_1
X_07010_ _07063_/A VGND VGND VPWR VPWR _07040_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08961_ _08962_/A _08962_/B VGND VGND VPWR VPWR _08966_/A sky130_fd_sc_hd__nor2_1
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07912_ _07912_/A _07912_/B VGND VGND VPWR VPWR _07916_/B sky130_fd_sc_hd__or2_1
X_08892_ _08867_/Y _08890_/Y _08987_/S VGND VGND VPWR VPWR _08893_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07843_ _07856_/B _07842_/X _07843_/S VGND VGND VPWR VPWR _07844_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07774_ _07786_/A _07786_/B VGND VGND VPWR VPWR _07783_/A sky130_fd_sc_hd__xnor2_1
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09513_ _09513_/A _09513_/B VGND VGND VPWR VPWR _09534_/A sky130_fd_sc_hd__nand2_1
X_06725_ _06725_/A VGND VGND VPWR VPWR _06727_/A sky130_fd_sc_hd__clkinv_2
XFILLER_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_157_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _14656_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09444_ _09437_/X _09442_/X _09443_/Y _08615_/X VGND VGND VPWR VPWR _13600_/D sky130_fd_sc_hd__a31o_1
X_06656_ _07804_/B _07804_/C VGND VGND VPWR VPWR _06656_/X sky130_fd_sc_hd__and2_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06587_ _12895_/Q _06580_/X _06586_/Y VGND VGND VPWR VPWR _12895_/D sky130_fd_sc_hd__o21a_1
X_09375_ _13591_/Q _09383_/B VGND VGND VPWR VPWR _09377_/B sky130_fd_sc_hd__or2_1
XFILLER_149_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08326_ _08340_/C VGND VGND VPWR VPWR _08331_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08257_ _08257_/A _08257_/B VGND VGND VPWR VPWR _08257_/Y sky130_fd_sc_hd__xnor2_1
X_07208_ _07208_/A _07208_/B VGND VGND VPWR VPWR _07209_/B sky130_fd_sc_hd__xnor2_1
Xclkbuf_3_5_0_clk clkbuf_3_5_0_clk/A VGND VGND VPWR VPWR clkbuf_3_5_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08188_ _13360_/Q _08188_/B VGND VGND VPWR VPWR _08189_/B sky130_fd_sc_hd__nor2_1
XFILLER_118_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07139_ _07139_/A _07190_/D VGND VGND VPWR VPWR _07147_/A sky130_fd_sc_hd__nand2_1
XFILLER_161_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10150_ _10150_/A _10150_/B VGND VGND VPWR VPWR _10150_/X sky130_fd_sc_hd__or2_1
XFILLER_106_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10081_ _10016_/A _10068_/X _10072_/X VGND VGND VPWR VPWR _10081_/X sky130_fd_sc_hd__a21o_1
XFILLER_87_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13840_ _14724_/CLK _13840_/D VGND VGND VPWR VPWR _13840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_148_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _14717_/CLK sky130_fd_sc_hd__clkbuf_16
X_13771_ _14720_/CLK _13771_/D VGND VGND VPWR VPWR _13771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10983_ _12645_/A _10980_/X _10982_/X _10929_/X VGND VGND VPWR VPWR _10983_/X sky130_fd_sc_hd__o211a_1
XFILLER_43_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12722_ _13606_/CLK _12722_/D VGND VGND VPWR VPWR hold454/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12653_ _14082_/CLK hold511/X _12609_/A VGND VGND VPWR VPWR hold496/A sky130_fd_sc_hd__dfrtp_1
XFILLER_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11604_ _13979_/Q _11446_/X _11612_/S VGND VGND VPWR VPWR _11605_/A sky130_fd_sc_hd__mux2_1
X_12584_ _12584_/A _14731_/Q VGND VGND VPWR VPWR _12584_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14323_ _14688_/CLK _14323_/D VGND VGND VPWR VPWR _14323_/Q sky130_fd_sc_hd__dfxtp_1
X_11535_ _13627_/Q _11541_/B VGND VGND VPWR VPWR _11536_/A sky130_fd_sc_hd__and2_1
XFILLER_128_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14254_ _14256_/CLK _14254_/D VGND VGND VPWR VPWR _14254_/Q sky130_fd_sc_hd__dfxtp_1
X_11466_ _11498_/A VGND VGND VPWR VPWR _11479_/S sky130_fd_sc_hd__buf_2
XFILLER_99_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13205_ _13604_/CLK _13205_/D VGND VGND VPWR VPWR hold80/A sky130_fd_sc_hd__dfxtp_1
X_10417_ _10418_/B _10417_/B VGND VGND VPWR VPWR _10426_/A sky130_fd_sc_hd__and2b_1
XFILLER_152_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14185_ _14201_/CLK _14185_/D VGND VGND VPWR VPWR _14185_/Q sky130_fd_sc_hd__dfxtp_1
X_11397_ _13722_/Q _11405_/B VGND VGND VPWR VPWR _11398_/A sky130_fd_sc_hd__and2_1
XFILLER_136_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13136_ _13359_/CLK _13136_/D hold1/X VGND VGND VPWR VPWR _13136_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _14624_/Q _10348_/B VGND VGND VPWR VPWR _13121_/D sky130_fd_sc_hd__xnor2_4
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10279_ _14325_/Q _14323_/Q _10593_/A VGND VGND VPWR VPWR _10279_/X sky130_fd_sc_hd__mux2_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _14555_/CLK _13067_/D VGND VGND VPWR VPWR hold392/A sky130_fd_sc_hd__dfxtp_1
X_12018_ _12018_/A VGND VGND VPWR VPWR _14315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_139_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _14159_/CLK sky130_fd_sc_hd__clkbuf_16
X_13969_ _13978_/CLK _13969_/D VGND VGND VPWR VPWR _13969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06510_ _06510_/A VGND VGND VPWR VPWR _12885_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07490_ _13149_/Q _09212_/B VGND VGND VPWR VPWR _07491_/B sky130_fd_sc_hd__or2_1
XFILLER_34_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06441_ _06455_/A _06532_/B _06444_/A VGND VGND VPWR VPWR _06446_/B sky130_fd_sc_hd__a21o_1
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09160_ _09161_/C _09160_/B _09146_/X VGND VGND VPWR VPWR _09160_/X sky130_fd_sc_hd__or3b_1
XFILLER_21_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06372_ hold479/X _10293_/A _14638_/D _06371_/X VGND VGND VPWR VPWR _13389_/D sky130_fd_sc_hd__a31o_1
XFILLER_147_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08111_ _08220_/B _08119_/C VGND VGND VPWR VPWR _08113_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09091_ _07570_/X _09089_/X _09090_/Y _07261_/X VGND VGND VPWR VPWR _13524_/D sky130_fd_sc_hd__a31o_1
XFILLER_148_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08042_ _10803_/A VGND VGND VPWR VPWR _08051_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_147_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09993_ _14647_/Q VGND VGND VPWR VPWR _10636_/A sky130_fd_sc_hd__clkbuf_2
X_08944_ _08944_/A _08944_/B VGND VGND VPWR VPWR _08944_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_131_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08875_ _08875_/A _08902_/B VGND VGND VPWR VPWR _08894_/B sky130_fd_sc_hd__nor2_1
XFILLER_56_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07826_ _13256_/Q _07832_/B VGND VGND VPWR VPWR _07833_/B sky130_fd_sc_hd__xnor2_1
XFILLER_29_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07757_ _07731_/A _07757_/B VGND VGND VPWR VPWR _07757_/X sky130_fd_sc_hd__and2b_1
XFILLER_72_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06708_ _06786_/A _06716_/A VGND VGND VPWR VPWR _06710_/B sky130_fd_sc_hd__xnor2_2
X_07688_ _07688_/A _07688_/B VGND VGND VPWR VPWR _07705_/A sky130_fd_sc_hd__nand2_1
XFILLER_52_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09427_ _09421_/A _09421_/B _09447_/A VGND VGND VPWR VPWR _09427_/X sky130_fd_sc_hd__o21ba_1
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06639_ _13032_/Q VGND VGND VPWR VPWR _07802_/A sky130_fd_sc_hd__buf_2
X_09358_ _09358_/A VGND VGND VPWR VPWR _12804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08309_ _08309_/A _08309_/B VGND VGND VPWR VPWR _13374_/D sky130_fd_sc_hd__nor2_1
XFILLER_139_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09289_ _13554_/Q _09289_/B VGND VGND VPWR VPWR _09289_/Y sky130_fd_sc_hd__xnor2_1
X_11320_ _14517_/Q VGND VGND VPWR VPWR _11320_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11251_ _11262_/A _11251_/B VGND VGND VPWR VPWR _11251_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10202_ _14398_/Q _14390_/Q _10627_/A VGND VGND VPWR VPWR _10626_/D sky130_fd_sc_hd__mux2_1
X_11182_ _14030_/Q _13996_/Q _13836_/Q _14548_/Q _11152_/X _11153_/X VGND VGND VPWR
+ VPWR _11183_/A sky130_fd_sc_hd__mux4_1
XFILLER_133_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10133_ _13867_/Q _13851_/Q _10137_/S VGND VGND VPWR VPWR _10134_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10064_ _14041_/D _10063_/X _14050_/D VGND VGND VPWR VPWR _10064_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13823_ _14533_/CLK _13823_/D VGND VGND VPWR VPWR _13823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13754_ _14644_/CLK _13754_/D VGND VGND VPWR VPWR _13754_/Q sky130_fd_sc_hd__dfxtp_1
X_10966_ _10966_/A _10925_/X VGND VGND VPWR VPWR _10966_/X sky130_fd_sc_hd__or2b_1
X_12705_ _13314_/CLK _12705_/D VGND VGND VPWR VPWR hold416/A sky130_fd_sc_hd__dfxtp_1
X_13685_ _13704_/CLK _13685_/D repeater56/X VGND VGND VPWR VPWR _13685_/Q sky130_fd_sc_hd__dfrtp_1
X_10897_ _14746_/Q _14736_/Q VGND VGND VPWR VPWR _10899_/C sky130_fd_sc_hd__xor2_1
XFILLER_70_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12636_ _14743_/Q _12635_/B _12609_/X VGND VGND VPWR VPWR _12637_/B sky130_fd_sc_hd__o21ai_1
XFILLER_34_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12567_ _12625_/B VGND VGND VPWR VPWR _12567_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14306_ _14543_/CLK _14306_/D VGND VGND VPWR VPWR _14306_/Q sky130_fd_sc_hd__dfxtp_1
X_11518_ _11518_/A VGND VGND VPWR VPWR _13840_/D sky130_fd_sc_hd__clkbuf_1
X_12498_ _12502_/A _12502_/B input16/X VGND VGND VPWR VPWR _12499_/A sky130_fd_sc_hd__and3_1
XFILLER_145_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold208 hold208/A VGND VGND VPWR VPWR hold208/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold219 hold219/A VGND VGND VPWR VPWR hold219/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_14237_ _14667_/CLK _14237_/D VGND VGND VPWR VPWR _14237_/Q sky130_fd_sc_hd__dfxtp_1
X_11449_ _11498_/A VGND VGND VPWR VPWR _11523_/S sky130_fd_sc_hd__buf_2
XFILLER_153_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14168_ _14209_/CLK hold326/X VGND VGND VPWR VPWR _14168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _13524_/CLK _13119_/D VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__dfxtp_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ _13027_/Q _08008_/B VGND VGND VPWR VPWR _06990_/Y sky130_fd_sc_hd__nand2_1
X_14099_ _14319_/CLK _14099_/D VGND VGND VPWR VPWR _14099_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05941_ _13875_/Q _13876_/Q _13877_/Q VGND VGND VPWR VPWR _05944_/A sky130_fd_sc_hd__or3_1
XFILLER_79_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08660_ _13450_/Q _09472_/B VGND VGND VPWR VPWR _08662_/A sky130_fd_sc_hd__and2_1
XFILLER_54_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07611_ _13112_/Q VGND VGND VPWR VPWR _07668_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08591_ _08591_/A VGND VGND VPWR VPWR _09424_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07542_ _13155_/Q _09289_/B _07548_/A _07547_/A VGND VGND VPWR VPWR _07543_/B sky130_fd_sc_hd__a22o_1
XFILLER_53_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07473_ _07473_/A _07586_/B VGND VGND VPWR VPWR _09215_/A sky130_fd_sc_hd__and2_1
X_09212_ _13542_/Q _09212_/B VGND VGND VPWR VPWR _09220_/D sky130_fd_sc_hd__xnor2_1
XFILLER_50_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06424_ _06500_/A _06421_/X _06422_/Y _06423_/Y VGND VGND VPWR VPWR _12878_/D sky130_fd_sc_hd__o31ai_1
X_06355_ _14686_/Q VGND VGND VPWR VPWR _06355_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_147_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09143_ _09161_/B _09161_/C _09141_/Y _09084_/A VGND VGND VPWR VPWR _09143_/X sky130_fd_sc_hd__o31a_1
XFILLER_148_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09074_ _09074_/A VGND VGND VPWR VPWR _12770_/D sky130_fd_sc_hd__clkbuf_1
X_06286_ _13953_/D _13954_/D _13955_/D _13956_/D VGND VGND VPWR VPWR _06287_/D sky130_fd_sc_hd__and4_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08025_ _08097_/A VGND VGND VPWR VPWR _10818_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_151_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09976_ _13754_/Q VGND VGND VPWR VPWR _10597_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08927_ _08927_/A _08978_/D VGND VGND VPWR VPWR _08935_/A sky130_fd_sc_hd__nand2_1
XFILLER_58_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08858_ _08870_/A _08870_/B VGND VGND VPWR VPWR _08860_/B sky130_fd_sc_hd__xnor2_1
XFILLER_73_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07809_ _06656_/X _07808_/X _07843_/S VGND VGND VPWR VPWR _07810_/A sky130_fd_sc_hd__mux2_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08789_ _08789_/A _08789_/B VGND VGND VPWR VPWR _08791_/A sky130_fd_sc_hd__nand2_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _10820_/A _13030_/Q VGND VGND VPWR VPWR _10821_/A sky130_fd_sc_hd__and2_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10751_ _12998_/Q _10820_/A VGND VGND VPWR VPWR _10752_/A sky130_fd_sc_hd__and2_1
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13470_ _13621_/CLK _13470_/D VGND VGND VPWR VPWR _13470_/Q sky130_fd_sc_hd__dfxtp_1
X_10682_ _10682_/A VGND VGND VPWR VPWR _12920_/D sky130_fd_sc_hd__clkbuf_1
X_14759__70 VGND VGND VPWR VPWR _14759__70/HI _13470_/D sky130_fd_sc_hd__conb_1
X_12421_ _12502_/B VGND VGND VPWR VPWR _12484_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_139_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12352_ _12352_/A VGND VGND VPWR VPWR _14599_/D sky130_fd_sc_hd__clkbuf_1
X_11303_ _11303_/A VGND VGND VPWR VPWR _13761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12283_ _14558_/Q _11950_/X _12291_/S VGND VGND VPWR VPWR _12284_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14022_ _14709_/CLK _14022_/D VGND VGND VPWR VPWR _14022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11234_ _14034_/Q _14000_/Q _13840_/Q _14552_/Q _10993_/A _10995_/A VGND VGND VPWR
+ VPWR _11235_/A sky130_fd_sc_hd__mux4_1
X_11165_ _11177_/A _11165_/B VGND VGND VPWR VPWR _11165_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10116_ _14185_/Q _14177_/Q _10617_/A VGND VGND VPWR VPWR _10116_/X sky130_fd_sc_hd__mux2_1
X_11096_ _11088_/X _11090_/Y _11094_/Y _11095_/X VGND VGND VPWR VPWR _11097_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10047_ _10047_/A VGND VGND VPWR VPWR _13949_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold80 hold80/A VGND VGND VPWR VPWR hold80/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold91 hold91/A VGND VGND VPWR VPWR hold91/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_90_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13806_ _13843_/CLK _13806_/D VGND VGND VPWR VPWR _13806_/Q sky130_fd_sc_hd__dfxtp_1
X_11998_ _14309_/Q _11997_/X _11998_/S VGND VGND VPWR VPWR _11999_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13737_ _13843_/CLK hold158/X VGND VGND VPWR VPWR _13737_/Q sky130_fd_sc_hd__dfxtp_1
X_10949_ _13318_/Q _10907_/X _10930_/X _10948_/Y VGND VGND VPWR VPWR _13318_/D sky130_fd_sc_hd__o22a_1
XFILLER_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_70_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _13423_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13668_ _14251_/CLK _13668_/D repeater56/X VGND VGND VPWR VPWR _13668_/Q sky130_fd_sc_hd__dfrtp_1
X_12619_ _12619_/A _12619_/B VGND VGND VPWR VPWR _12619_/X sky130_fd_sc_hd__or2_1
XFILLER_129_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13599_ _13621_/CLK _13599_/D repeater56/X VGND VGND VPWR VPWR _13599_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06140_ _14188_/Q _14180_/Q _14194_/D VGND VGND VPWR VPWR _06145_/C sky130_fd_sc_hd__mux2_1
XFILLER_145_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_0 _12025_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06071_ _13957_/Q _13949_/Q _13962_/D VGND VGND VPWR VPWR _06075_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09830_ _09830_/A _09830_/B VGND VGND VPWR VPWR _09840_/A sky130_fd_sc_hd__or2_1
XFILLER_99_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _09761_/A _09761_/B VGND VGND VPWR VPWR _09763_/A sky130_fd_sc_hd__or2_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ _06981_/A _06973_/B _06973_/C VGND VGND VPWR VPWR _06973_/Y sky130_fd_sc_hd__nand3_1
XFILLER_39_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _13455_/Q _09511_/B VGND VGND VPWR VPWR _08713_/B sky130_fd_sc_hd__or2_1
X_05924_ _13843_/D _13713_/Q _13714_/Q _13715_/Q VGND VGND VPWR VPWR _05924_/X sky130_fd_sc_hd__and4_1
XFILLER_100_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09692_ _09720_/A _09709_/C VGND VGND VPWR VPWR _09695_/B sky130_fd_sc_hd__and2_1
XFILLER_39_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08643_ _08633_/X _08641_/Y _08642_/X VGND VGND VPWR VPWR _13448_/D sky130_fd_sc_hd__a21o_1
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08574_ _08622_/A _08574_/B VGND VGND VPWR VPWR _08590_/B sky130_fd_sc_hd__or2_1
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07525_ _07515_/A _07519_/X _07532_/C _07524_/X VGND VGND VPWR VPWR _07525_/X sky130_fd_sc_hd__a31o_1
XFILLER_41_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_61_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _14636_/CLK sky130_fd_sc_hd__clkbuf_16
X_07456_ _07411_/X _07453_/X _07454_/Y _07455_/X VGND VGND VPWR VPWR _13146_/D sky130_fd_sc_hd__a31o_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06407_ _06401_/X _06402_/Y _06405_/X _06586_/A VGND VGND VPWR VPWR _12877_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_109_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07387_ _07387_/A VGND VGND VPWR VPWR _07400_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_157_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09126_ _13530_/Q _09126_/B VGND VGND VPWR VPWR _09134_/D sky130_fd_sc_hd__xnor2_1
XFILLER_148_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06338_ _06338_/A VGND VGND VPWR VPWR _14404_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06269_ _13807_/Q _13791_/Q _06281_/S VGND VGND VPWR VPWR _06270_/A sky130_fd_sc_hd__mux2_1
X_09057_ _09057_/A VGND VGND VPWR VPWR _12762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08008_ _13281_/Q _08008_/B VGND VGND VPWR VPWR _08008_/X sky130_fd_sc_hd__or2_1
XFILLER_150_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09959_ _13700_/Q VGND VGND VPWR VPWR _09968_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_58_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12970_ _12970_/CLK hold321/X VGND VGND VPWR VPWR _12970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11921_ _14267_/Q _11481_/X _11929_/S VGND VGND VPWR VPWR _11922_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _14644_/CLK _14640_/D VGND VGND VPWR VPWR _14640_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _11852_/A VGND VGND VPWR VPWR _14224_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10803_ _10803_/A VGND VGND VPWR VPWR _10812_/B sky130_fd_sc_hd__clkbuf_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _14605_/CLK _14571_/D VGND VGND VPWR VPWR _14571_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _11783_/A VGND VGND VPWR VPWR _14085_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_52_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _14647_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13522_ _13596_/CLK _13522_/D VGND VGND VPWR VPWR _13522_/Q sky130_fd_sc_hd__dfxtp_1
X_10734_ _12901_/Q _10742_/B VGND VGND VPWR VPWR _10735_/A sky130_fd_sc_hd__and2_1
XFILLER_158_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13453_ _13605_/CLK _13453_/D repeater57/X VGND VGND VPWR VPWR _13453_/Q sky130_fd_sc_hd__dfrtp_1
X_10665_ _10665_/A _10665_/B VGND VGND VPWR VPWR _12914_/D sky130_fd_sc_hd__nor2_1
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12404_ _10596_/B _12404_/B VGND VGND VPWR VPWR _12405_/A sky130_fd_sc_hd__and2b_1
XFILLER_127_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13384_ _14530_/CLK _13384_/D _12609_/A VGND VGND VPWR VPWR _13384_/Q sky130_fd_sc_hd__dfrtp_1
X_10596_ _14629_/Q _10596_/B VGND VGND VPWR VPWR _14621_/D sky130_fd_sc_hd__xor2_1
XFILLER_154_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12335_ _12335_/A VGND VGND VPWR VPWR _14591_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12266_ _11343_/X _14548_/Q _12270_/S VGND VGND VPWR VPWR _12267_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14005_ _14679_/CLK _14005_/D VGND VGND VPWR VPWR _14005_/Q sky130_fd_sc_hd__dfxtp_1
X_11217_ _11240_/A _11217_/B VGND VGND VPWR VPWR _11217_/Y sky130_fd_sc_hd__nor2_1
X_12197_ _12197_/A VGND VGND VPWR VPWR _14509_/D sky130_fd_sc_hd__clkbuf_1
X_11148_ _11179_/A _11148_/B VGND VGND VPWR VPWR _11148_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11079_ _12645_/B VGND VGND VPWR VPWR _11079_/X sky130_fd_sc_hd__buf_2
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_43_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _12881_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07310_ _09099_/A _07302_/B _07311_/C _07461_/A VGND VGND VPWR VPWR _07313_/A sky130_fd_sc_hd__a22o_1
X_08290_ _08301_/C VGND VGND VPWR VPWR _08294_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07241_ _07241_/A VGND VGND VPWR VPWR _07311_/A sky130_fd_sc_hd__clkbuf_2
X_07172_ _07139_/A _07203_/B _07147_/B _07171_/X VGND VGND VPWR VPWR _07174_/B sky130_fd_sc_hd__a31oi_2
XFILLER_158_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06123_ _06122_/X _06116_/X _06127_/A VGND VGND VPWR VPWR _06124_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06054_ _06054_/A VGND VGND VPWR VPWR _13917_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09813_ _09813_/A VGND VGND VPWR VPWR _09816_/A sky130_fd_sc_hd__inv_2
XFILLER_100_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09744_ _09673_/X _09685_/X _09688_/X _09718_/Y VGND VGND VPWR VPWR _09746_/B sky130_fd_sc_hd__o22a_1
X_06956_ _06968_/A _06967_/A VGND VGND VPWR VPWR _06956_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05907_ _13807_/Q _13808_/Q _13809_/Q _13810_/Q VGND VGND VPWR VPWR _05909_/B sky130_fd_sc_hd__and4_1
X_09675_ _09715_/S _14213_/Q VGND VGND VPWR VPWR _09675_/X sky130_fd_sc_hd__or2b_1
X_06887_ _06887_/A _06887_/B VGND VGND VPWR VPWR _06924_/A sky130_fd_sc_hd__nand2_1
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08626_ _08657_/A _08624_/X _08634_/A VGND VGND VPWR VPWR _09451_/B sky130_fd_sc_hd__o21a_1
XFILLER_55_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _13442_/Q _09407_/B _09407_/C VGND VGND VPWR VPWR _08572_/B sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_34_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _12974_/CLK sky130_fd_sc_hd__clkbuf_16
X_07508_ _07477_/B _07505_/Y _07507_/X VGND VGND VPWR VPWR _07510_/B sky130_fd_sc_hd__a21oi_1
X_08488_ _14250_/Q _14246_/Q _14248_/Q _13712_/Q _08473_/C _08545_/S VGND VGND VPWR
+ VPWR _08488_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07439_ _07400_/A _07330_/X _07435_/A VGND VGND VPWR VPWR _07444_/A sky130_fd_sc_hd__o21a_2
XFILLER_155_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10450_ _10450_/A _10468_/A VGND VGND VPWR VPWR _10452_/A sky130_fd_sc_hd__or2_1
XFILLER_10_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09109_ _09109_/A _09109_/B _09109_/C VGND VGND VPWR VPWR _09134_/A sky130_fd_sc_hd__or3_1
X_10381_ _13516_/Q _13519_/Q _13520_/Q _14211_/D VGND VGND VPWR VPWR _10387_/B sky130_fd_sc_hd__a22o_1
XFILLER_108_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12120_ _14475_/Q _11984_/X _12128_/S VGND VGND VPWR VPWR _12121_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12051_ _12051_/A VGND VGND VPWR VPWR _14444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold380 hold380/A VGND VGND VPWR VPWR hold380/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold391 hold391/A VGND VGND VPWR VPWR hold391/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11002_ _14261_/Q _14652_/Q _13759_/Q _14707_/Q _10940_/X _10942_/X VGND VGND VPWR
+ VPWR _11003_/B sky130_fd_sc_hd__mux4_1
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12953_ _13039_/CLK hold293/X VGND VGND VPWR VPWR _12953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11904_ _11904_/A VGND VGND VPWR VPWR _14259_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12884_ _12885_/CLK _12884_/D hold1/X VGND VGND VPWR VPWR _12884_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _14636_/CLK _14623_/D VGND VGND VPWR VPWR _14623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11835_ _11835_/A VGND VGND VPWR VPWR _14109_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _13574_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14725_/CLK _14554_/D VGND VGND VPWR VPWR _14554_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _11375_/X _14074_/Q _11766_/S VGND VGND VPWR VPWR _11767_/A sky130_fd_sc_hd__mux2_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13505_ _13855_/CLK hold274/X VGND VGND VPWR VPWR _13505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10717_ _10717_/A VGND VGND VPWR VPWR _12936_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14485_ _14617_/CLK _14485_/D VGND VGND VPWR VPWR _14485_/Q sky130_fd_sc_hd__dfxtp_1
X_11697_ _11697_/A VGND VGND VPWR VPWR _14030_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13436_ _14010_/CLK _13436_/D repeater56/X VGND VGND VPWR VPWR _13436_/Q sky130_fd_sc_hd__dfrtp_1
X_10648_ _10648_/A VGND VGND VPWR VPWR _12672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13367_ _13423_/CLK _13367_/D repeater56/X VGND VGND VPWR VPWR _13367_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10579_ hold159/A hold59/A VGND VGND VPWR VPWR _10580_/A sky130_fd_sc_hd__or2_1
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12318_ _14574_/Q _12004_/X _12324_/S VGND VGND VPWR VPWR _12319_/A sky130_fd_sc_hd__mux2_1
X_13298_ _13298_/CLK hold440/X VGND VGND VPWR VPWR _13298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12249_ _12249_/A VGND VGND VPWR VPWR _14540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06810_ _13008_/Q _07876_/B VGND VGND VPWR VPWR _06820_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07790_ _07790_/A _07790_/B VGND VGND VPWR VPWR _07791_/B sky130_fd_sc_hd__xnor2_1
XFILLER_84_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06741_ _06895_/A VGND VGND VPWR VPWR _06743_/A sky130_fd_sc_hd__clkbuf_4
X_09460_ _09460_/A _09460_/B VGND VGND VPWR VPWR _09466_/B sky130_fd_sc_hd__and2_1
X_06672_ _13346_/Q _13344_/Q _06705_/S VGND VGND VPWR VPWR _06672_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08411_ _08411_/A VGND VGND VPWR VPWR _12736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09391_ _09391_/A _09391_/B _09390_/X VGND VGND VPWR VPWR _09419_/A sky130_fd_sc_hd__or3b_2
Xclkbuf_leaf_16_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _14413_/CLK sky130_fd_sc_hd__clkbuf_16
X_08342_ _08340_/X _09084_/A _08342_/C VGND VGND VPWR VPWR _08343_/A sky130_fd_sc_hd__and3b_1
XFILLER_60_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08273_ _08273_/A _08273_/B VGND VGND VPWR VPWR _08283_/A sky130_fd_sc_hd__or2_1
X_07224_ _07224_/A VGND VGND VPWR VPWR _07461_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_164_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07155_ _07155_/A _07182_/B VGND VGND VPWR VPWR _07156_/B sky130_fd_sc_hd__nand2_1
XFILLER_106_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06106_ _06106_/A VGND VGND VPWR VPWR _13943_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07086_ _07083_/Y _07114_/A _07086_/C _13707_/Q VGND VGND VPWR VPWR _07114_/B sky130_fd_sc_hd__and4bb_1
XFILLER_161_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06037_ hold42/A _10293_/A VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__nand2_2
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07988_ _13278_/Q _07988_/B VGND VGND VPWR VPWR _07995_/A sky130_fd_sc_hd__nand2_1
XFILLER_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09727_ _13701_/Q VGND VGND VPWR VPWR _09855_/A sky130_fd_sc_hd__clkbuf_2
X_06939_ _13020_/Q _06954_/A VGND VGND VPWR VPWR _06940_/B sky130_fd_sc_hd__nor2_1
XFILLER_16_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09658_ _09720_/A VGND VGND VPWR VPWR _09758_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ _08591_/A _08607_/B _08607_/C _08596_/A VGND VGND VPWR VPWR _09440_/C sky130_fd_sc_hd__o22ai_4
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _09600_/A VGND VGND VPWR VPWR _09598_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11620_ _11620_/A VGND VGND VPWR VPWR _13986_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11551_ _11551_/A VGND VGND VPWR VPWR _13858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10502_ _10502_/A VGND VGND VPWR VPWR _14012_/D sky130_fd_sc_hd__clkbuf_1
X_14270_ _14716_/CLK _14270_/D VGND VGND VPWR VPWR _14270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11482_ _11498_/A VGND VGND VPWR VPWR _11495_/S sky130_fd_sc_hd__buf_2
XFILLER_137_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13221_ _13423_/CLK hold453/X VGND VGND VPWR VPWR _13221_/Q sky130_fd_sc_hd__dfxtp_1
X_10433_ hold71/A VGND VGND VPWR VPWR _10485_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13152_ _13372_/CLK _13152_/D repeater57/X VGND VGND VPWR VPWR _13152_/Q sky130_fd_sc_hd__dfrtp_1
X_10364_ _10415_/A _10376_/A VGND VGND VPWR VPWR _10366_/B sky130_fd_sc_hd__or2_1
XFILLER_3_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12103_ _12103_/A VGND VGND VPWR VPWR _14467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _13528_/CLK hold289/X VGND VGND VPWR VPWR _13083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10295_ _10601_/A _10296_/B _10601_/C VGND VGND VPWR VPWR _13816_/D sky130_fd_sc_hd__nand3_1
XFILLER_105_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12034_ _14684_/Q _12034_/B VGND VGND VPWR VPWR _12035_/A sky130_fd_sc_hd__and2_1
XFILLER_78_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13985_ _14539_/CLK _13985_/D VGND VGND VPWR VPWR _13985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12936_ _12970_/CLK _12936_/D VGND VGND VPWR VPWR hold133/A sky130_fd_sc_hd__dfxtp_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12867_ _13811_/CLK _12867_/D VGND VGND VPWR VPWR hold346/A sky130_fd_sc_hd__dfxtp_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14606_ _14714_/CLK _14606_/D VGND VGND VPWR VPWR _14606_/Q sky130_fd_sc_hd__dfxtp_1
X_11818_ _11818_/A VGND VGND VPWR VPWR _14101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12798_ _13570_/CLK _12798_/D VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__dfxtp_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _14737_/CLK _14537_/D VGND VGND VPWR VPWR _14537_/Q sky130_fd_sc_hd__dfxtp_1
X_11749_ _11749_/A VGND VGND VPWR VPWR _11758_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_14_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14468_ _14705_/CLK _14468_/D VGND VGND VPWR VPWR _14468_/Q sky130_fd_sc_hd__dfxtp_1
X_13419_ _14696_/CLK hold85/X VGND VGND VPWR VPWR _13419_/Q sky130_fd_sc_hd__dfxtp_1
X_14399_ _14732_/CLK _14399_/D VGND VGND VPWR VPWR _14399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08960_ _08927_/A _08991_/B _08935_/B _08959_/X VGND VGND VPWR VPWR _08962_/B sky130_fd_sc_hd__a31oi_1
Xclkbuf_leaf_5_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _14275_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07911_ _13267_/Q _07911_/B VGND VGND VPWR VPWR _07912_/B sky130_fd_sc_hd__nor2_1
X_08891_ _09006_/S VGND VGND VPWR VPWR _08987_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_96_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07842_ _07858_/C _07842_/B VGND VGND VPWR VPWR _07842_/X sky130_fd_sc_hd__xor2_1
XFILLER_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07773_ _07773_/A _07773_/B VGND VGND VPWR VPWR _07786_/B sky130_fd_sc_hd__nor2_1
XFILLER_83_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09512_ _13609_/Q _09518_/B VGND VGND VPWR VPWR _09513_/B sky130_fd_sc_hd__or2_1
XFILLER_25_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06724_ _13003_/Q _07840_/B VGND VGND VPWR VPWR _06725_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09443_ _09443_/A _09443_/B _09454_/D VGND VGND VPWR VPWR _09443_/Y sky130_fd_sc_hd__nand3_1
X_06655_ _06881_/B _06652_/C _06652_/D _06881_/A VGND VGND VPWR VPWR _07804_/C sky130_fd_sc_hd__a22o_1
XFILLER_13_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09374_ _13589_/Q _09370_/B _09368_/X _09369_/A VGND VGND VPWR VPWR _09377_/A sky130_fd_sc_hd__a31o_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06586_ _06586_/A _06595_/B VGND VGND VPWR VPWR _06586_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08325_ _13378_/Q _13379_/Q _13380_/Q _08325_/D VGND VGND VPWR VPWR _08340_/C sky130_fd_sc_hd__and4_1
XFILLER_149_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08256_ _08256_/A _08256_/B VGND VGND VPWR VPWR _08257_/B sky130_fd_sc_hd__nand2_1
XFILLER_137_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07207_ _07207_/A _07207_/B VGND VGND VPWR VPWR _07208_/B sky130_fd_sc_hd__xnor2_1
X_08187_ _13360_/Q _08188_/B VGND VGND VPWR VPWR _08189_/A sky130_fd_sc_hd__and2_1
XFILLER_152_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07138_ _07138_/A VGND VGND VPWR VPWR _13347_/D sky130_fd_sc_hd__clkbuf_1
X_07069_ _07069_/A _07069_/B VGND VGND VPWR VPWR _07082_/B sky130_fd_sc_hd__xnor2_1
XFILLER_79_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10080_ _10080_/A VGND VGND VPWR VPWR _13902_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13770_ _14667_/CLK _13770_/D VGND VGND VPWR VPWR _13770_/Q sky130_fd_sc_hd__dfxtp_1
X_10982_ _10982_/A _10925_/X VGND VGND VPWR VPWR _10982_/X sky130_fd_sc_hd__or2b_1
XFILLER_55_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12721_ _13604_/CLK _12721_/D VGND VGND VPWR VPWR hold342/A sky130_fd_sc_hd__dfxtp_1
XFILLER_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12652_ _14082_/CLK hold175/X _12609_/A VGND VGND VPWR VPWR hold511/A sky130_fd_sc_hd__dfrtp_1
XFILLER_90_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11603_ _11653_/S VGND VGND VPWR VPWR _11612_/S sky130_fd_sc_hd__buf_2
X_12583_ _14746_/Q _14731_/Q VGND VGND VPWR VPWR _12583_/X sky130_fd_sc_hd__or2_1
XFILLER_156_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14322_ _14425_/CLK hold281/X VGND VGND VPWR VPWR hold117/A sky130_fd_sc_hd__dfxtp_1
X_11534_ _11534_/A VGND VGND VPWR VPWR _13850_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14253_ _14256_/CLK _14253_/D VGND VGND VPWR VPWR _14253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11465_ _14699_/Q VGND VGND VPWR VPWR _11465_/X sky130_fd_sc_hd__clkbuf_2
X_13204_ _13606_/CLK _13204_/D VGND VGND VPWR VPWR hold517/A sky130_fd_sc_hd__dfxtp_1
X_10416_ _10416_/A _10416_/B VGND VGND VPWR VPWR _10417_/B sky130_fd_sc_hd__nor2_1
XFILLER_143_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14184_ _14196_/CLK _14184_/D VGND VGND VPWR VPWR _14184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11396_ _11444_/B VGND VGND VPWR VPWR _11405_/B sky130_fd_sc_hd__clkbuf_1
X_13135_ _13534_/CLK _13135_/D hold1/X VGND VGND VPWR VPWR _13135_/Q sky130_fd_sc_hd__dfrtp_1
X_10347_ _10347_/A _10347_/B VGND VGND VPWR VPWR _13038_/D sky130_fd_sc_hd__xnor2_1
XFILLER_152_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _14082_/CLK _13066_/D VGND VGND VPWR VPWR hold451/A sky130_fd_sc_hd__dfxtp_1
X_10278_ _10278_/A VGND VGND VPWR VPWR _12663_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12017_ _14315_/Q _12016_/X _12026_/S VGND VGND VPWR VPWR _12018_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13968_ _13978_/CLK _13968_/D VGND VGND VPWR VPWR _13968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12919_ _13039_/CLK _12919_/D VGND VGND VPWR VPWR hold235/A sky130_fd_sc_hd__dfxtp_1
X_13899_ _14693_/CLK hold273/X VGND VGND VPWR VPWR hold95/A sky130_fd_sc_hd__dfxtp_1
X_06440_ _14439_/Q _14437_/Q _06458_/S VGND VGND VPWR VPWR _06532_/B sky130_fd_sc_hd__mux2_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06371_ _06044_/B _06371_/B input22/X VGND VGND VPWR VPWR _06371_/X sky130_fd_sc_hd__and3b_1
XFILLER_148_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08110_ _08208_/A _08209_/B _08108_/X _08147_/A VGND VGND VPWR VPWR _08119_/C sky130_fd_sc_hd__a22o_1
X_09090_ _09089_/A _09089_/B _09089_/C VGND VGND VPWR VPWR _09090_/Y sky130_fd_sc_hd__o21ai_1
X_08041_ _08041_/A VGND VGND VPWR VPWR _12682_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09992_ _09992_/A VGND VGND VPWR VPWR _13708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08943_ _08943_/A _08970_/B VGND VGND VPWR VPWR _08944_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_15_0_clk clkbuf_3_7_0_clk/X VGND VGND VPWR VPWR clkbuf_4_15_0_clk/X sky130_fd_sc_hd__clkbuf_2
X_08874_ _08871_/Y _08902_/A _08874_/C _13518_/D VGND VGND VPWR VPWR _08902_/B sky130_fd_sc_hd__and4bb_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07825_ _07825_/A VGND VGND VPWR VPWR _13255_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07756_ _07756_/A _07756_/B VGND VGND VPWR VPWR _07760_/B sky130_fd_sc_hd__and2_1
XFILLER_71_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06707_ _06881_/A _06720_/B VGND VGND VPWR VPWR _06716_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07687_ _07687_/A VGND VGND VPWR VPWR _13659_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09426_ _09447_/D VGND VGND VPWR VPWR _09454_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06638_ _06881_/B _06652_/C VGND VGND VPWR VPWR _07807_/B sky130_fd_sc_hd__xor2_4
XFILLER_13_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09357_ _13314_/Q _13552_/Q _10822_/A VGND VGND VPWR VPWR _09358_/A sky130_fd_sc_hd__mux2_1
X_06569_ _06569_/A _06569_/B VGND VGND VPWR VPWR _06569_/Y sky130_fd_sc_hd__xnor2_1
X_08308_ _13374_/Q _08314_/B _08338_/A VGND VGND VPWR VPWR _08309_/B sky130_fd_sc_hd__o21ai_1
X_09288_ _08218_/X _09286_/X _09287_/Y _07526_/X VGND VGND VPWR VPWR _13553_/D sky130_fd_sc_hd__a31o_1
XFILLER_21_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08239_ _08232_/B _08237_/Y _08286_/S VGND VGND VPWR VPWR _08240_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11250_ _14279_/Q _14670_/Q _13777_/Q _14725_/Q _10914_/A _10918_/A VGND VGND VPWR
+ VPWR _11251_/B sky130_fd_sc_hd__mux4_1
XFILLER_107_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10201_ _10201_/A VGND VGND VPWR VPWR _14417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11181_ _14312_/Q _14482_/Q _14238_/Q _14068_/Q _11137_/X _11138_/X VGND VGND VPWR
+ VPWR _11181_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10132_ _10132_/A VGND VGND VPWR VPWR _14180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10063_ _10063_/A _10063_/B VGND VGND VPWR VPWR _10063_/X sky130_fd_sc_hd__or2_1
XFILLER_85_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13822_ _14533_/CLK _13822_/D VGND VGND VPWR VPWR _13822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13753_ _14633_/CLK _13753_/D VGND VGND VPWR VPWR hold208/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10965_ _14015_/Q _13981_/Q _13821_/Q _14533_/Q _10921_/X _10922_/X VGND VGND VPWR
+ VPWR _10966_/A sky130_fd_sc_hd__mux4_1
XFILLER_62_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12704_ _13314_/CLK _12704_/D VGND VGND VPWR VPWR hold76/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13684_ _13686_/CLK _13684_/D repeater56/X VGND VGND VPWR VPWR _13684_/Q sky130_fd_sc_hd__dfrtp_1
X_10896_ _14745_/Q _14735_/Q VGND VGND VPWR VPWR _10899_/B sky130_fd_sc_hd__xor2_1
XFILLER_31_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12635_ _14743_/Q _12635_/B VGND VGND VPWR VPWR _12637_/A sky130_fd_sc_hd__and2_1
XFILLER_31_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12566_ _12566_/A VGND VGND VPWR VPWR _12625_/B sky130_fd_sc_hd__inv_2
XFILLER_8_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14305_ _14602_/CLK _14305_/D VGND VGND VPWR VPWR _14305_/Q sky130_fd_sc_hd__dfxtp_1
X_11517_ _13840_/Q _11516_/X _11523_/S VGND VGND VPWR VPWR _11518_/A sky130_fd_sc_hd__mux2_1
X_12497_ _12497_/A VGND VGND VPWR VPWR _14678_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14236_ _14667_/CLK _14236_/D VGND VGND VPWR VPWR _14236_/Q sky130_fd_sc_hd__dfxtp_1
Xhold209 hold209/A VGND VGND VPWR VPWR hold209/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_11448_ _12150_/A _12226_/A VGND VGND VPWR VPWR _11498_/A sky130_fd_sc_hd__nor2_8
XFILLER_109_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14167_ _14209_/CLK _14167_/D VGND VGND VPWR VPWR hold326/A sky130_fd_sc_hd__dfxtp_1
X_11379_ _11379_/A VGND VGND VPWR VPWR _13783_/D sky130_fd_sc_hd__clkbuf_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _14679_/CLK hold131/X VGND VGND VPWR VPWR hold394/A sky130_fd_sc_hd__dfxtp_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14098_ _14098_/CLK _14098_/D VGND VGND VPWR VPWR _14098_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05940_ hold199/A _13862_/Q _13863_/Q _13866_/Q VGND VGND VPWR VPWR _05945_/C sky130_fd_sc_hd__or4_1
XFILLER_85_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13049_ _13528_/CLK _13049_/D VGND VGND VPWR VPWR hold343/A sky130_fd_sc_hd__dfxtp_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07610_ _07610_/A _07610_/B VGND VGND VPWR VPWR _07614_/A sky130_fd_sc_hd__nor2_1
XFILLER_94_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08590_ _08590_/A _08590_/B _08622_/B VGND VGND VPWR VPWR _08590_/X sky130_fd_sc_hd__and3_1
Xclkbuf_3_4_0_clk clkbuf_3_5_0_clk/A VGND VGND VPWR VPWR clkbuf_4_9_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07541_ _07586_/B VGND VGND VPWR VPWR _09289_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_81_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07472_ _07579_/B VGND VGND VPWR VPWR _07586_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_09211_ _09182_/X _09214_/B _09210_/Y _07575_/X VGND VGND VPWR VPWR _13541_/D sky130_fd_sc_hd__a31o_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06423_ _06586_/A _06423_/B VGND VGND VPWR VPWR _06423_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09142_ _09161_/B _09161_/C _09141_/Y VGND VGND VPWR VPWR _09142_/Y sky130_fd_sc_hd__o21ai_1
X_06354_ _14685_/Q _12034_/B _14590_/D _14681_/Q VGND VGND VPWR VPWR _12874_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09073_ _13234_/Q _13463_/Q _09075_/S VGND VGND VPWR VPWR _09074_/A sky130_fd_sc_hd__mux2_1
X_06285_ _13957_/D _13958_/D _13959_/D VGND VGND VPWR VPWR _06287_/C sky130_fd_sc_hd__and3_1
XFILLER_136_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08024_ hold23/A VGND VGND VPWR VPWR _08097_/A sky130_fd_sc_hd__buf_2
XFILLER_162_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09975_ _09975_/A VGND VGND VPWR VPWR _12873_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08926_ _08926_/A VGND VGND VPWR VPWR _14250_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08857_ _08857_/A _08857_/B VGND VGND VPWR VPWR _08870_/B sky130_fd_sc_hd__xnor2_1
XFILLER_58_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07808_ _07808_/A _07808_/B VGND VGND VPWR VPWR _07808_/X sky130_fd_sc_hd__xor2_1
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08788_ _13465_/Q _09576_/B VGND VGND VPWR VPWR _08789_/B sky130_fd_sc_hd__or2_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07739_ _07718_/Y _07738_/Y _07781_/S VGND VGND VPWR VPWR _07740_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10750_ _10781_/A VGND VGND VPWR VPWR _10820_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09409_ _13595_/Q _09417_/B VGND VGND VPWR VPWR _09409_/Y sky130_fd_sc_hd__nand2_1
X_10681_ _12877_/Q _10687_/B VGND VGND VPWR VPWR _10682_/A sky130_fd_sc_hd__and2_1
XFILLER_41_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12420_ _12502_/A VGND VGND VPWR VPWR _12484_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_127_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12351_ _14599_/Q _11962_/X _12353_/S VGND VGND VPWR VPWR _12352_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11302_ _13761_/Q _11301_/X _11311_/S VGND VGND VPWR VPWR _11303_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12282_ _12332_/S VGND VGND VPWR VPWR _12291_/S sky130_fd_sc_hd__buf_2
XFILLER_4_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14021_ _14697_/CLK _14021_/D VGND VGND VPWR VPWR _14021_/Q sky130_fd_sc_hd__dfxtp_1
X_11233_ _14316_/Q _14486_/Q _14242_/Q _14072_/Q _11208_/X _11209_/X VGND VGND VPWR
+ VPWR _11233_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11164_ _14272_/Q _14663_/Q _13770_/Q _14718_/Q _11162_/X _11163_/X VGND VGND VPWR
+ VPWR _11165_/B sky130_fd_sc_hd__mux4_1
XFILLER_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10115_ _14181_/Q _14173_/Q _10617_/A VGND VGND VPWR VPWR _10616_/D sky130_fd_sc_hd__mux2_1
X_11095_ _11166_/A VGND VGND VPWR VPWR _11095_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10046_ _13803_/Q _13787_/Q _10050_/S VGND VGND VPWR VPWR _10047_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold70 hold70/A VGND VGND VPWR VPWR hold70/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold81 hold81/A VGND VGND VPWR VPWR hold81/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold92 hold92/A VGND VGND VPWR VPWR hold92/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_64_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13805_ _13805_/CLK _13805_/D VGND VGND VPWR VPWR _13805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11997_ _14519_/Q VGND VGND VPWR VPWR _11997_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10948_ _10948_/A _12626_/B VGND VGND VPWR VPWR _10948_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13736_ _13805_/CLK hold130/X VGND VGND VPWR VPWR _13736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10879_ _13156_/Q _10885_/B VGND VGND VPWR VPWR _10880_/A sky130_fd_sc_hd__and2_1
X_13667_ _14251_/CLK _13667_/D repeater56/X VGND VGND VPWR VPWR _13667_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12618_ _11655_/A _12619_/B _12616_/X _12617_/X VGND VGND VPWR VPWR _14736_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13598_ _13598_/CLK _13598_/D repeater56/X VGND VGND VPWR VPWR _13598_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_129_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12549_ _12549_/A VGND VGND VPWR VPWR _14719_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1 _11636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06070_ _13956_/Q _13948_/Q _13962_/D VGND VGND VPWR VPWR _06075_/C sky130_fd_sc_hd__mux2_1
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14219_ _14440_/CLK _14219_/D VGND VGND VPWR VPWR _14219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09760_ _13674_/Q _09760_/B VGND VGND VPWR VPWR _09761_/B sky130_fd_sc_hd__nor2_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06972_ _06973_/B _06973_/C _06981_/A VGND VGND VPWR VPWR _06978_/B sky130_fd_sc_hd__a21o_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _13455_/Q _08746_/A VGND VGND VPWR VPWR _08713_/A sky130_fd_sc_hd__nand2_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05923_ _13716_/Q _13717_/Q _13718_/Q _13719_/Q VGND VGND VPWR VPWR _05923_/X sky130_fd_sc_hd__and4_1
X_09691_ _09685_/X _09827_/B _09687_/X _09688_/X _09787_/S _09736_/A VGND VGND VPWR
+ VPWR _09709_/C sky130_fd_sc_hd__mux4_1
XFILLER_67_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08642_ _08642_/A _09457_/B _09457_/C VGND VGND VPWR VPWR _08642_/X sky130_fd_sc_hd__and3_1
XFILLER_55_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08573_ _08539_/X _08572_/Y _08558_/A VGND VGND VPWR VPWR _08574_/B sky130_fd_sc_hd__a21o_1
XFILLER_19_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07524_ _08157_/A VGND VGND VPWR VPWR _07524_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_35_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07455_ _07455_/A _09188_/B VGND VGND VPWR VPWR _07455_/X sky130_fd_sc_hd__and2_1
XFILLER_22_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06406_ _06500_/A VGND VGND VPWR VPWR _06586_/A sky130_fd_sc_hd__buf_2
XFILLER_10_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07386_ _07327_/X _07461_/B _07461_/A VGND VGND VPWR VPWR _07389_/A sky130_fd_sc_hd__o21ai_2
X_09125_ _09125_/A VGND VGND VPWR VPWR _09125_/X sky130_fd_sc_hd__buf_2
XFILLER_157_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06337_ _14105_/Q _14089_/Q _10224_/S VGND VGND VPWR VPWR _06338_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09056_ _13226_/Q _13455_/Q _09064_/S VGND VGND VPWR VPWR _09057_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06268_ _06273_/S VGND VGND VPWR VPWR _06281_/S sky130_fd_sc_hd__clkbuf_2
X_08007_ _13281_/Q _08008_/B VGND VGND VPWR VPWR _08007_/Y sky130_fd_sc_hd__nand2_1
XFILLER_150_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06199_ _06199_/A VGND VGND VPWR VPWR _14367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09958_ _09958_/A VGND VGND VPWR VPWR _12865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08909_ _08909_/A _08909_/B VGND VGND VPWR VPWR _08911_/C sky130_fd_sc_hd__xnor2_1
X_09889_ _13695_/Q _09893_/A _09894_/A VGND VGND VPWR VPWR _09889_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11920_ _11931_/A VGND VGND VPWR VPWR _11929_/S sky130_fd_sc_hd__buf_2
XFILLER_73_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _14224_/Q _11459_/X _11853_/S VGND VGND VPWR VPWR _11852_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _10802_/A VGND VGND VPWR VPWR _13063_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _14610_/CLK _14570_/D VGND VGND VPWR VPWR _14570_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11782_ _13563_/Q _11784_/B VGND VGND VPWR VPWR _11783_/A sky130_fd_sc_hd__and2_1
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10733_ _13031_/D VGND VGND VPWR VPWR _10742_/B sky130_fd_sc_hd__clkbuf_1
X_13521_ _13704_/CLK hold504/X VGND VGND VPWR VPWR hold207/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13452_ _13602_/CLK _13452_/D repeater57/X VGND VGND VPWR VPWR _13452_/Q sky130_fd_sc_hd__dfrtp_1
X_10664_ _14339_/Q _10666_/C _10656_/X VGND VGND VPWR VPWR _10665_/B sky130_fd_sc_hd__o21ai_1
XFILLER_13_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12403_ _12403_/A VGND VGND VPWR VPWR _14628_/D sky130_fd_sc_hd__clkbuf_1
X_13383_ _14333_/CLK _13383_/D _12609_/A VGND VGND VPWR VPWR _13383_/Q sky130_fd_sc_hd__dfrtp_1
X_10595_ _13699_/Q _13704_/Q hold508/X _09776_/X VGND VGND VPWR VPWR _13699_/D sky130_fd_sc_hd__o31a_1
XFILLER_139_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12334_ _14639_/Q _12340_/B _12336_/C VGND VGND VPWR VPWR _12335_/A sky130_fd_sc_hd__and3_1
XFILLER_56_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12265_ _12265_/A VGND VGND VPWR VPWR _14547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14004_ _14679_/CLK _14004_/D VGND VGND VPWR VPWR _14004_/Q sky130_fd_sc_hd__dfxtp_1
X_11216_ _14276_/Q _14667_/Q _13774_/Q _14722_/Q _11162_/X _11163_/X VGND VGND VPWR
+ VPWR _11217_/B sky130_fd_sc_hd__mux4_1
X_12196_ _14509_/Q _12016_/X _12202_/S VGND VGND VPWR VPWR _12197_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11147_ _11088_/X _11144_/Y _11146_/Y _11095_/X VGND VGND VPWR VPWR _11148_/B sky130_fd_sc_hd__a211o_1
XFILLER_68_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11078_ _13327_/Q _11008_/X _11071_/X _11077_/Y VGND VGND VPWR VPWR _13327_/D sky130_fd_sc_hd__o22a_1
XFILLER_95_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10029_ _13953_/Q _13945_/Q _10607_/A VGND VGND VPWR VPWR _10029_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13719_ _13799_/CLK hold179/X VGND VGND VPWR VPWR _13719_/Q sky130_fd_sc_hd__dfxtp_1
X_14699_ _14710_/CLK hold306/X VGND VGND VPWR VPWR _14699_/Q sky130_fd_sc_hd__dfxtp_1
X_07240_ _13167_/Q VGND VGND VPWR VPWR _07241_/A sky130_fd_sc_hd__inv_2
XFILLER_31_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07171_ _07146_/B _07171_/B VGND VGND VPWR VPWR _07171_/X sky130_fd_sc_hd__and2b_1
XFILLER_9_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06122_ _14202_/Q _14200_/Q _14209_/Q VGND VGND VPWR VPWR _06122_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06053_ _06052_/X _06046_/X _06057_/A VGND VGND VPWR VPWR _06054_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09812_ _09812_/A _09812_/B VGND VGND VPWR VPWR _09813_/A sky130_fd_sc_hd__or2_1
XFILLER_113_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06955_ _13022_/Q _07981_/B VGND VGND VPWR VPWR _06967_/A sky130_fd_sc_hd__xor2_1
X_09743_ _09743_/A VGND VGND VPWR VPWR _13672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05906_ _13811_/Q _13812_/Q _13813_/Q VGND VGND VPWR VPWR _05909_/A sky130_fd_sc_hd__and3_1
XFILLER_28_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09674_ _09688_/S VGND VGND VPWR VPWR _09715_/S sky130_fd_sc_hd__clkbuf_2
X_06886_ _13014_/Q _07947_/B VGND VGND VPWR VPWR _06887_/B sky130_fd_sc_hd__or2_1
XFILLER_39_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _09424_/B _08596_/B _08607_/C _08566_/B VGND VGND VPWR VPWR _08634_/A sky130_fd_sc_hd__o31a_1
XFILLER_43_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08556_ _13442_/Q _08556_/B VGND VGND VPWR VPWR _08558_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07507_ _13147_/Q _13148_/Q _13149_/Q _13150_/Q _09257_/B VGND VGND VPWR VPWR _07507_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_51_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08487_ _13473_/Q _14254_/Q _14256_/Q _14252_/Q _08473_/C _08545_/S VGND VGND VPWR
+ VPWR _08606_/B sky130_fd_sc_hd__mux4_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07438_ _07438_/A _07438_/B VGND VGND VPWR VPWR _07443_/A sky130_fd_sc_hd__nor2_1
XFILLER_149_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07369_ _07416_/A _07369_/B VGND VGND VPWR VPWR _07369_/X sky130_fd_sc_hd__or2_1
X_09108_ _09095_/A _09095_/B _09101_/Y _09099_/X VGND VGND VPWR VPWR _09109_/C sky130_fd_sc_hd__o211a_1
XFILLER_164_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10380_ _10398_/B _10380_/B VGND VGND VPWR VPWR _14215_/D sky130_fd_sc_hd__xnor2_1
XFILLER_164_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09039_ _09039_/A VGND VGND VPWR VPWR _12755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12050_ _11291_/X _14444_/Q _12052_/S VGND VGND VPWR VPWR _12051_/A sky130_fd_sc_hd__mux2_1
Xhold370 hold370/A VGND VGND VPWR VPWR hold370/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_105_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold381 hold381/A VGND VGND VPWR VPWR hold381/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_11001_ _11001_/A VGND VGND VPWR VPWR _11001_/Y sky130_fd_sc_hd__inv_2
Xhold392 hold392/A VGND VGND VPWR VPWR hold392/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12952_ _13039_/CLK hold235/X VGND VGND VPWR VPWR _12952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11903_ _14259_/Q _11456_/X _11907_/S VGND VGND VPWR VPWR _11904_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _12930_/CLK _12883_/D hold1/X VGND VGND VPWR VPWR _12883_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _14645_/CLK _14622_/D VGND VGND VPWR VPWR _14622_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_93_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ hold173/A _11834_/B VGND VGND VPWR VPWR _11835_/A sky130_fd_sc_hd__and2_1
XFILLER_73_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _11765_/A VGND VGND VPWR VPWR _14073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14553_ _14725_/CLK _14553_/D VGND VGND VPWR VPWR _14553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _13855_/CLK hold435/X VGND VGND VPWR VPWR _13504_/Q sky130_fd_sc_hd__dfxtp_1
X_10716_ _12893_/Q _10720_/B VGND VGND VPWR VPWR _10717_/A sky130_fd_sc_hd__and2_1
X_14484_ _14510_/CLK _14484_/D VGND VGND VPWR VPWR _14484_/Q sky130_fd_sc_hd__dfxtp_1
X_11696_ _14030_/Q _11504_/X _11700_/S VGND VGND VPWR VPWR _11697_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10647_ _10647_/A _10647_/B VGND VGND VPWR VPWR _10648_/A sky130_fd_sc_hd__and2_1
X_13435_ _13476_/CLK _13435_/D repeater56/X VGND VGND VPWR VPWR _13435_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_155_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13366_ _13366_/CLK _13366_/D repeater56/X VGND VGND VPWR VPWR _13366_/Q sky130_fd_sc_hd__dfrtp_1
X_10578_ hold159/A _12911_/Q _12908_/Q _06542_/X VGND VGND VPWR VPWR _12908_/D sky130_fd_sc_hd__o31a_1
X_12317_ _12317_/A VGND VGND VPWR VPWR _14573_/D sky130_fd_sc_hd__clkbuf_1
X_13297_ _13303_/CLK hold389/X VGND VGND VPWR VPWR _13297_/Q sky130_fd_sc_hd__dfxtp_1
X_12248_ _11310_/X _14540_/Q _12248_/S VGND VGND VPWR VPWR _12249_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12179_ _14501_/Q _11991_/X _12183_/S VGND VGND VPWR VPWR _12180_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06740_ _06730_/A _06730_/B _06725_/A _06727_/B _06739_/Y VGND VGND VPWR VPWR _06740_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_92_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06671_ _06671_/A VGND VGND VPWR VPWR _06852_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08410_ _13100_/Q _08331_/A _08418_/S VGND VGND VPWR VPWR _08411_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09390_ _13592_/Q _08495_/B _09377_/A _09377_/B _09383_/X VGND VGND VPWR VPWR _09390_/X
+ sky130_fd_sc_hd__a221o_1
X_08341_ _08331_/A _08331_/B _08340_/D _13384_/Q VGND VGND VPWR VPWR _08342_/C sky130_fd_sc_hd__a31o_1
XFILLER_32_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08272_ _13368_/Q _08272_/B VGND VGND VPWR VPWR _08273_/B sky130_fd_sc_hd__nor2_1
XFILLER_149_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07223_ _13169_/Q VGND VGND VPWR VPWR _07224_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07154_ _07153_/A _07153_/B _07153_/C VGND VGND VPWR VPWR _07182_/B sky130_fd_sc_hd__o21ai_2
XFILLER_146_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06105_ _13797_/Q _06105_/B VGND VGND VPWR VPWR _06106_/A sky130_fd_sc_hd__and2_1
XFILLER_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07085_ _07086_/C _13707_/Q _07083_/Y _07114_/A VGND VGND VPWR VPWR _07087_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_106_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06036_ _06371_/B VGND VGND VPWR VPWR _10293_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07987_ _07987_/A _07987_/B VGND VGND VPWR VPWR _07992_/C sky130_fd_sc_hd__nand2_1
XFILLER_86_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06938_ _13020_/Q _06938_/B VGND VGND VPWR VPWR _06948_/A sky130_fd_sc_hd__and2_1
X_09726_ _09726_/A _09726_/B VGND VGND VPWR VPWR _09726_/X sky130_fd_sc_hd__xor2_1
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06869_ _06870_/A _06870_/B _06876_/B VGND VGND VPWR VPWR _06869_/X sky130_fd_sc_hd__a21o_1
X_09657_ _13703_/Q VGND VGND VPWR VPWR _09720_/A sky130_fd_sc_hd__inv_2
XFILLER_103_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _08671_/C VGND VGND VPWR VPWR _09440_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09588_ _09588_/A VGND VGND VPWR VPWR _12809_/D sky130_fd_sc_hd__buf_2
XFILLER_42_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _08530_/A _08530_/B _08525_/A _08527_/B _08538_/Y VGND VGND VPWR VPWR _08539_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11550_ _13634_/Q _11552_/B VGND VGND VPWR VPWR _11551_/A sky130_fd_sc_hd__and2_1
XFILLER_23_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10501_ _10485_/C _10503_/B _10501_/C VGND VGND VPWR VPWR _10502_/A sky130_fd_sc_hd__and3b_1
XFILLER_11_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11481_ _14515_/Q VGND VGND VPWR VPWR _11481_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13220_ _13606_/CLK hold348/X VGND VGND VPWR VPWR _13220_/Q sky130_fd_sc_hd__dfxtp_1
X_10432_ _10432_/A _10432_/B VGND VGND VPWR VPWR _14212_/D sky130_fd_sc_hd__nor2_1
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13151_ _13555_/CLK _13151_/D repeater57/X VGND VGND VPWR VPWR _13151_/Q sky130_fd_sc_hd__dfrtp_1
X_10363_ _13516_/Q VGND VGND VPWR VPWR _10376_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12102_ _14467_/Q _11959_/X _12106_/S VGND VGND VPWR VPWR _12103_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13082_ _13528_/CLK hold343/X VGND VGND VPWR VPWR _13082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10294_ input1/X input12/X _12402_/B VGND VGND VPWR VPWR _10601_/C sky130_fd_sc_hd__o21ai_1
XFILLER_3_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12033_ _12033_/A VGND VGND VPWR VPWR _14325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13984_ _14536_/CLK _13984_/D VGND VGND VPWR VPWR _13984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12935_ _12970_/CLK _12935_/D VGND VGND VPWR VPWR hold359/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _13811_/CLK _12866_/D VGND VGND VPWR VPWR hold172/A sky130_fd_sc_hd__dfxtp_1
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _14605_/CLK _14605_/D VGND VGND VPWR VPWR _14605_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11817_ _13579_/Q _11817_/B VGND VGND VPWR VPWR _11818_/A sky130_fd_sc_hd__and2_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _13570_/CLK _12797_/D VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__dfxtp_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ _14536_/CLK _14536_/D VGND VGND VPWR VPWR _14536_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11748_ _11748_/A VGND VGND VPWR VPWR _14065_/D sky130_fd_sc_hd__clkbuf_1
X_14467_ _14742_/CLK _14467_/D VGND VGND VPWR VPWR _14467_/Q sky130_fd_sc_hd__dfxtp_1
X_11679_ _11679_/A VGND VGND VPWR VPWR _14022_/D sky130_fd_sc_hd__clkbuf_1
X_13418_ _13617_/CLK hold104/X VGND VGND VPWR VPWR _13418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14398_ _14410_/CLK _14398_/D VGND VGND VPWR VPWR _14398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13349_ _14432_/CLK _13349_/D VGND VGND VPWR VPWR _13349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07910_ _13267_/Q _07910_/B VGND VGND VPWR VPWR _07912_/A sky130_fd_sc_hd__and2_1
XFILLER_130_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08890_ _08944_/A _08890_/B VGND VGND VPWR VPWR _08890_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_123_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07841_ _07835_/A _07858_/A _07839_/Y _07840_/Y VGND VGND VPWR VPWR _07842_/B sky130_fd_sc_hd__a31o_1
XFILLER_68_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07772_ _07772_/A _07772_/B _07785_/C _07772_/D VGND VGND VPWR VPWR _07773_/B sky130_fd_sc_hd__and4_1
XFILLER_83_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09511_ _13609_/Q _09511_/B VGND VGND VPWR VPWR _09513_/A sky130_fd_sc_hd__nand2_1
X_06723_ _06723_/A VGND VGND VPWR VPWR _07840_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_52_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09442_ _09443_/A _09443_/B _09454_/D VGND VGND VPWR VPWR _09442_/X sky130_fd_sc_hd__a21o_1
X_06654_ _06736_/A VGND VGND VPWR VPWR _06881_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09373_ _09373_/A VGND VGND VPWR VPWR _13590_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06585_ _06598_/C VGND VGND VPWR VPWR _06595_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08324_ _13379_/Q _08322_/A _08323_/Y VGND VGND VPWR VPWR _13379_/D sky130_fd_sc_hd__a21oi_1
XFILLER_33_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08255_ _08236_/A _08245_/Y _08236_/B _08244_/A _08233_/A VGND VGND VPWR VPWR _08256_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_20_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07206_ _07206_/A _07206_/B VGND VGND VPWR VPWR _07207_/B sky130_fd_sc_hd__nor2_1
X_08186_ _08199_/A _08186_/B _08186_/C VGND VGND VPWR VPWR _08188_/B sky130_fd_sc_hd__and3_1
XFILLER_118_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07137_ _07102_/Y _07136_/Y _07199_/S VGND VGND VPWR VPWR _07138_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07068_ _14634_/Q hold154/A VGND VGND VPWR VPWR _07069_/B sky130_fd_sc_hd__nand2_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06019_ _13558_/Q _06019_/B VGND VGND VPWR VPWR _06019_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09709_ _09778_/B _13669_/Q _09709_/C VGND VGND VPWR VPWR _09709_/X sky130_fd_sc_hd__and3_1
X_10981_ _14016_/Q _13982_/Q _13822_/Q _14534_/Q _10921_/X _10922_/X VGND VGND VPWR
+ VPWR _10982_/A sky130_fd_sc_hd__mux4_1
XFILLER_83_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12720_ _13596_/CLK _12720_/D VGND VGND VPWR VPWR hold463/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12651_ _13587_/CLK _13700_/D _12609_/A VGND VGND VPWR VPWR hold175/A sky130_fd_sc_hd__dfrtp_1
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11602_ _11636_/A VGND VGND VPWR VPWR _11653_/S sky130_fd_sc_hd__buf_2
XFILLER_70_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12582_ _12582_/A VGND VGND VPWR VPWR _12616_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14321_ _14536_/CLK hold117/X VGND VGND VPWR VPWR hold114/A sky130_fd_sc_hd__dfxtp_1
XFILLER_7_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11533_ _13626_/Q _11541_/B VGND VGND VPWR VPWR _11534_/A sky130_fd_sc_hd__and2_1
XFILLER_156_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14252_ _14256_/CLK _14252_/D VGND VGND VPWR VPWR _14252_/Q sky130_fd_sc_hd__dfxtp_1
X_11464_ _11464_/A VGND VGND VPWR VPWR _13823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10415_ _10415_/A _10429_/C _10415_/C VGND VGND VPWR VPWR _10416_/B sky130_fd_sc_hd__and3_1
X_13203_ _13372_/CLK _13203_/D VGND VGND VPWR VPWR hold201/A sky130_fd_sc_hd__dfxtp_1
X_14183_ _14209_/CLK _14183_/D VGND VGND VPWR VPWR _14183_/Q sky130_fd_sc_hd__dfxtp_1
X_11395_ _11395_/A VGND VGND VPWR VPWR _13790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13134_ _13534_/CLK _13134_/D hold1/X VGND VGND VPWR VPWR _13134_/Q sky130_fd_sc_hd__dfrtp_1
X_10346_ _10346_/A _13120_/D VGND VGND VPWR VPWR _10347_/B sky130_fd_sc_hd__xnor2_1
XFILLER_125_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _14082_/CLK _13065_/D VGND VGND VPWR VPWR hold372/A sky130_fd_sc_hd__dfxtp_1
X_10277_ _10272_/X _12508_/B _10592_/B VGND VGND VPWR VPWR _10278_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12016_ _12016_/A VGND VGND VPWR VPWR _12016_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13967_ _13978_/CLK _13967_/D VGND VGND VPWR VPWR _13967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12918_ _14710_/CLK _12918_/D VGND VGND VPWR VPWR hold384/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13898_ _14693_/CLK hold331/X VGND VGND VPWR VPWR hold339/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _13721_/CLK _12849_/D VGND VGND VPWR VPWR hold200/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06370_ hold473/X _10293_/A _14638_/D _06369_/X VGND VGND VPWR VPWR _13388_/D sky130_fd_sc_hd__a31o_1
XFILLER_9_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14519_ _14608_/CLK _14519_/D VGND VGND VPWR VPWR _14519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08040_ _12958_/Q _13258_/Q _08040_/S VGND VGND VPWR VPWR _08041_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09991_ _09990_/X _09987_/X _09991_/S VGND VGND VPWR VPWR _09992_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08942_ _08941_/A _08941_/B _08941_/C VGND VGND VPWR VPWR _08970_/B sky130_fd_sc_hd__o21ai_2
XFILLER_130_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08873_ _08874_/C _13518_/D _08871_/Y _08902_/A VGND VGND VPWR VPWR _08875_/A sky130_fd_sc_hd__o2bb2a_1
X_07824_ _07819_/B _07823_/Y _07843_/S VGND VGND VPWR VPWR _07825_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07755_ _07756_/A _07756_/B VGND VGND VPWR VPWR _07760_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06706_ _06630_/A _06704_/X _06705_/X _06633_/X _06674_/C _06745_/A VGND VGND VPWR
+ VPWR _06720_/B sky130_fd_sc_hd__mux4_1
X_07686_ _07661_/Y _07684_/Y _07781_/S VGND VGND VPWR VPWR _07687_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09425_ _09424_/B _09424_/C _13598_/Q VGND VGND VPWR VPWR _09447_/D sky130_fd_sc_hd__a21oi_1
X_06637_ _06671_/A _06633_/X _06634_/X _06767_/B _06636_/Y VGND VGND VPWR VPWR _06652_/C
+ sky130_fd_sc_hd__a32o_4
XFILLER_25_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09356_ _10831_/A VGND VGND VPWR VPWR _10822_/A sky130_fd_sc_hd__buf_4
X_06568_ _06567_/Y _06560_/B _06557_/A VGND VGND VPWR VPWR _06569_/B sky130_fd_sc_hd__a21oi_1
XFILLER_100_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08307_ _13374_/Q _08314_/B VGND VGND VPWR VPWR _08309_/A sky130_fd_sc_hd__and2_1
X_09287_ _09287_/A _09287_/B _09287_/C VGND VGND VPWR VPWR _09287_/Y sky130_fd_sc_hd__nand3_1
XFILLER_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06499_ _06499_/A _06499_/B _06499_/C VGND VGND VPWR VPWR _06499_/Y sky130_fd_sc_hd__nor3_1
X_08238_ _13165_/Q VGND VGND VPWR VPWR _08286_/S sky130_fd_sc_hd__buf_2
XFILLER_4_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08169_ _08169_/A _08169_/B VGND VGND VPWR VPWR _08170_/B sky130_fd_sc_hd__or2_1
XFILLER_107_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10200_ _10626_/C _10198_/X _10206_/S VGND VGND VPWR VPWR _10201_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11180_ _13334_/Q _11150_/X _11173_/X _11179_/Y VGND VGND VPWR VPWR _13334_/D sky130_fd_sc_hd__o22a_1
XFILLER_122_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10131_ _13866_/Q _13850_/Q _14167_/D VGND VGND VPWR VPWR _10132_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10062_ _14038_/D _10062_/B VGND VGND VPWR VPWR _10063_/B sky130_fd_sc_hd__nor2_1
XFILLER_48_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13821_ _14533_/CLK _13821_/D VGND VGND VPWR VPWR _13821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13752_ _14633_/CLK hold208/X VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__dfxtp_2
X_10964_ _14297_/Q _14467_/Q _14223_/Q _14053_/Q _10914_/X _12643_/A VGND VGND VPWR
+ VPWR _10964_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12703_ _13314_/CLK _12703_/D VGND VGND VPWR VPWR hold81/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13683_ _13686_/CLK _13683_/D repeater56/X VGND VGND VPWR VPWR _13683_/Q sky130_fd_sc_hd__dfrtp_1
X_10895_ _14748_/Q _14738_/Q VGND VGND VPWR VPWR _10899_/A sky130_fd_sc_hd__xor2_1
XFILLER_70_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12634_ _12634_/A VGND VGND VPWR VPWR _14742_/D sky130_fd_sc_hd__clkbuf_1
X_12565_ _12623_/B VGND VGND VPWR VPWR _12619_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14304_ _14495_/CLK _14304_/D VGND VGND VPWR VPWR _14304_/Q sky130_fd_sc_hd__dfxtp_1
X_11516_ _12019_/A VGND VGND VPWR VPWR _11516_/X sky130_fd_sc_hd__clkbuf_2
X_12496_ _12496_/A _12496_/B input15/X VGND VGND VPWR VPWR _12497_/A sky130_fd_sc_hd__and3_1
X_14235_ _14652_/CLK _14235_/D VGND VGND VPWR VPWR _14235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11447_ _12149_/A _11841_/A VGND VGND VPWR VPWR _12226_/A sky130_fd_sc_hd__nand2_8
XFILLER_4_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14166_ _14196_/CLK _14166_/D VGND VGND VPWR VPWR _14166_/Q sky130_fd_sc_hd__dfxtp_1
X_11378_ _13714_/Q _11382_/B VGND VGND VPWR VPWR _11379_/A sky130_fd_sc_hd__and2_1
XFILLER_113_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _13532_/CLK hold159/X VGND VGND VPWR VPWR hold507/A sky130_fd_sc_hd__dfxtp_1
X_10329_ _10329_/A _10329_/B VGND VGND VPWR VPWR _13171_/D sky130_fd_sc_hd__xnor2_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _14319_/CLK _14097_/D VGND VGND VPWR VPWR _14097_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _13528_/CLK _13048_/D VGND VGND VPWR VPWR hold121/A sky130_fd_sc_hd__dfxtp_1
XFILLER_112_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07540_ _13156_/Q _09257_/B VGND VGND VPWR VPWR _07547_/B sky130_fd_sc_hd__xor2_1
XFILLER_62_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07471_ _09277_/B VGND VGND VPWR VPWR _07579_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09210_ _09210_/A _09210_/B _09220_/C VGND VGND VPWR VPWR _09210_/Y sky130_fd_sc_hd__nand3_1
X_06422_ _06436_/A _06421_/C _06421_/A VGND VGND VPWR VPWR _06422_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09141_ _13531_/Q _07365_/X _09137_/Y VGND VGND VPWR VPWR _09141_/Y sky130_fd_sc_hd__a21oi_1
X_06353_ _06353_/A VGND VGND VPWR VPWR _12034_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_147_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09072_ _09072_/A VGND VGND VPWR VPWR _12769_/D sky130_fd_sc_hd__clkbuf_1
X_06284_ _13957_/D _13958_/D _13959_/D _06284_/D VGND VGND VPWR VPWR _06284_/X sky130_fd_sc_hd__or4_1
XFILLER_107_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08023_ _08021_/Y _08022_/X _07932_/A VGND VGND VPWR VPWR _13283_/D sky130_fd_sc_hd__o21bai_1
XFILLER_135_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09974_ _13510_/Q _13699_/Q _09974_/S VGND VGND VPWR VPWR _09975_/A sky130_fd_sc_hd__mux2_2
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08925_ _08890_/Y _08924_/Y _08987_/S VGND VGND VPWR VPWR _08926_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08856_ _13515_/D _13431_/Q VGND VGND VPWR VPWR _08857_/B sky130_fd_sc_hd__nand2_1
XFILLER_73_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07807_ _13252_/Q _07807_/B VGND VGND VPWR VPWR _07808_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05999_ _13565_/Q _13566_/Q _13567_/Q _13568_/Q VGND VGND VPWR VPWR _06002_/C sky130_fd_sc_hd__or4_1
X_08787_ _13465_/Q _08787_/B VGND VGND VPWR VPWR _08789_/A sky130_fd_sc_hd__nand2_1
XFILLER_85_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07738_ _07738_/A _07738_/B VGND VGND VPWR VPWR _07738_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07669_ _07669_/A _07696_/B VGND VGND VPWR VPWR _07688_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09408_ _09408_/A _09420_/A VGND VGND VPWR VPWR _09419_/D sky130_fd_sc_hd__or2_2
XFILLER_41_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10680_ _10680_/A VGND VGND VPWR VPWR _12919_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09339_ _13306_/Q _13544_/Q _09343_/S VGND VGND VPWR VPWR _09340_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12350_ _12350_/A VGND VGND VPWR VPWR _14598_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11301_ _14700_/Q VGND VGND VPWR VPWR _11301_/X sky130_fd_sc_hd__clkbuf_2
X_12281_ _12315_/A VGND VGND VPWR VPWR _12332_/S sky130_fd_sc_hd__buf_2
XFILLER_107_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11232_ _13338_/Q _10962_/A _11225_/X _11231_/Y VGND VGND VPWR VPWR _13338_/D sky130_fd_sc_hd__o22a_1
X_14020_ _14710_/CLK _14020_/D VGND VGND VPWR VPWR _14020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11163_ _11163_/A VGND VGND VPWR VPWR _11163_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10114_ _10114_/A VGND VGND VPWR VPWR _14200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11094_ _11106_/A _11094_/B VGND VGND VPWR VPWR _11094_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10045_ _10045_/A VGND VGND VPWR VPWR _13948_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold71 hold71/A VGND VGND VPWR VPWR hold71/X sky130_fd_sc_hd__clkbuf_2
Xhold82 hold82/A VGND VGND VPWR VPWR hold82/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold93 hold93/A VGND VGND VPWR VPWR hold93/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_91_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13804_ _13843_/CLK _13804_/D VGND VGND VPWR VPWR _13804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11996_ _11996_/A VGND VGND VPWR VPWR _14308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13735_ _13805_/CLK hold127/X VGND VGND VPWR VPWR _13735_/Q sky130_fd_sc_hd__dfxtp_1
X_10947_ _10932_/X _10938_/Y _10944_/Y _10946_/X VGND VGND VPWR VPWR _10948_/A sky130_fd_sc_hd__a211o_1
XFILLER_32_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13666_ _13666_/CLK _13666_/D VGND VGND VPWR VPWR _13666_/Q sky130_fd_sc_hd__dfxtp_1
X_10878_ _10878_/A VGND VGND VPWR VPWR _13197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12617_ _12641_/A VGND VGND VPWR VPWR _12617_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_14_0_clk clkbuf_3_7_0_clk/X VGND VGND VPWR VPWR clkbuf_4_14_0_clk/X sky130_fd_sc_hd__clkbuf_2
X_13597_ _13598_/CLK _13597_/D repeater56/X VGND VGND VPWR VPWR _13597_/Q sky130_fd_sc_hd__dfrtp_1
X_12548_ _11337_/X _14719_/Q _12554_/S VGND VGND VPWR VPWR _12549_/A sky130_fd_sc_hd__mux2_1
X_12479_ _12479_/A VGND VGND VPWR VPWR _14670_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_2 _11636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14218_ _14440_/CLK _14218_/D VGND VGND VPWR VPWR _14218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14149_ _14153_/CLK _14149_/D VGND VGND VPWR VPWR _14149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ _06978_/A _06971_/B VGND VGND VPWR VPWR _06981_/A sky130_fd_sc_hd__nand2_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _08706_/X _08708_/X _08709_/Y _08696_/X VGND VGND VPWR VPWR _13454_/D sky130_fd_sc_hd__a31o_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05922_ _13843_/D _13721_/Q _05915_/X _05917_/X _05921_/Y VGND VGND VPWR VPWR _05937_/A
+ sky130_fd_sc_hd__a41o_1
X_09690_ _13711_/Q VGND VGND VPWR VPWR _09736_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08641_ _08641_/A _08644_/B VGND VGND VPWR VPWR _08641_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_39_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08572_ _08572_/A _08572_/B VGND VGND VPWR VPWR _08572_/Y sky130_fd_sc_hd__nor2_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07523_ _07515_/A _07519_/X _07532_/C VGND VGND VPWR VPWR _07530_/B sky130_fd_sc_hd__a21oi_1
XFILLER_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07454_ _07454_/A _07454_/B _07454_/C VGND VGND VPWR VPWR _07454_/Y sky130_fd_sc_hd__nand3_1
XFILLER_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06405_ _10349_/A _06405_/B VGND VGND VPWR VPWR _06405_/X sky130_fd_sc_hd__and2_1
X_07385_ _07385_/A VGND VGND VPWR VPWR _13140_/D sky130_fd_sc_hd__clkbuf_1
X_06336_ _06336_/A VGND VGND VPWR VPWR _14403_/D sky130_fd_sc_hd__clkbuf_1
X_09124_ _08157_/X _07356_/B _09122_/X _09123_/Y VGND VGND VPWR VPWR _13529_/D sky130_fd_sc_hd__a22o_1
XFILLER_108_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09055_ _09600_/A VGND VGND VPWR VPWR _09064_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_135_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06267_ _06267_/A VGND VGND VPWR VPWR _13952_/D sky130_fd_sc_hd__clkbuf_1
X_08006_ _08004_/Y _08005_/X _07932_/A VGND VGND VPWR VPWR _13280_/D sky130_fd_sc_hd__o21bai_1
XFILLER_123_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06198_ _06196_/X _06192_/X _10193_/A VGND VGND VPWR VPWR _06199_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09957_ _13502_/Q _13691_/Q _09957_/S VGND VGND VPWR VPWR _09958_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08908_ _08908_/A _08938_/A VGND VGND VPWR VPWR _08909_/B sky130_fd_sc_hd__nor2_1
XFILLER_106_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _09893_/A _09888_/B VGND VGND VPWR VPWR _13694_/D sky130_fd_sc_hd__nor2_1
X_08839_ _08846_/B _08839_/B VGND VGND VPWR VPWR _08841_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _11850_/A VGND VGND VPWR VPWR _14223_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10801_ _13021_/Q _10801_/B VGND VGND VPWR VPWR _10802_/A sky130_fd_sc_hd__and2_1
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11781_ _11781_/A VGND VGND VPWR VPWR _14084_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13520_ _13520_/CLK _13520_/D VGND VGND VPWR VPWR _13520_/Q sky130_fd_sc_hd__dfxtp_1
X_10732_ _10732_/A VGND VGND VPWR VPWR _12943_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13451_ _13700_/CLK _13451_/D repeater57/X VGND VGND VPWR VPWR _13451_/Q sky130_fd_sc_hd__dfrtp_1
X_10663_ _14339_/Q _10666_/C VGND VGND VPWR VPWR _10665_/A sky130_fd_sc_hd__and2_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12402_ _06044_/B _12402_/B input20/X VGND VGND VPWR VPWR _12403_/A sky130_fd_sc_hd__and3b_1
X_10594_ _14583_/Q _14590_/Q VGND VGND VPWR VPWR _13748_/D sky130_fd_sc_hd__xor2_1
X_13382_ _14530_/CLK _13382_/D _12609_/A VGND VGND VPWR VPWR _13382_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12333_ _12333_/A VGND VGND VPWR VPWR _14581_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_clk clkbuf_3_3_0_clk/A VGND VGND VPWR VPWR clkbuf_4_7_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_126_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12264_ _11337_/X _14547_/Q _12270_/S VGND VGND VPWR VPWR _12265_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14003_ _14679_/CLK hold46/X VGND VGND VPWR VPWR _14003_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_107_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11215_ _11215_/A VGND VGND VPWR VPWR _11215_/Y sky130_fd_sc_hd__inv_2
X_12195_ _12195_/A VGND VGND VPWR VPWR _14508_/D sky130_fd_sc_hd__clkbuf_1
Xoutput50 _13324_/Q VGND VGND VPWR VPWR data_o[6] sky130_fd_sc_hd__buf_2
XFILLER_150_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11146_ _11177_/A _11146_/B VGND VGND VPWR VPWR _11146_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11077_ _11108_/A _11077_/B VGND VGND VPWR VPWR _11077_/Y sky130_fd_sc_hd__nand2_1
XFILLER_163_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10028_ _13949_/Q _13941_/Q _10607_/A VGND VGND VPWR VPWR _10606_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11979_ _14303_/Q _11978_/X _11982_/S VGND VGND VPWR VPWR _11980_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13718_ _13727_/CLK hold436/X VGND VGND VPWR VPWR _13718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14698_ _14710_/CLK hold102/X VGND VGND VPWR VPWR _14698_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13649_ _14327_/CLK hold312/X VGND VGND VPWR VPWR _13649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07170_ _07190_/D VGND VGND VPWR VPWR _07203_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06121_ _06121_/A VGND VGND VPWR VPWR _14148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_120_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _14180_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06052_ _13970_/Q _13968_/Q _13977_/Q VGND VGND VPWR VPWR _06052_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09811_ _13679_/Q _09811_/B VGND VGND VPWR VPWR _09812_/B sky130_fd_sc_hd__nor2_1
XFILLER_86_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09742_ _09739_/B _09741_/X _09774_/S VGND VGND VPWR VPWR _09743_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06954_ _06954_/A VGND VGND VPWR VPWR _07981_/B sky130_fd_sc_hd__buf_2
XFILLER_39_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05905_ hold52/A _13798_/Q _13799_/Q _13802_/Q VGND VGND VPWR VPWR _05910_/C sky130_fd_sc_hd__and4_1
X_09673_ _09718_/A _13711_/Q VGND VGND VPWR VPWR _09673_/X sky130_fd_sc_hd__or2b_1
Xclkbuf_leaf_187_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _14704_/CLK sky130_fd_sc_hd__clkbuf_16
X_06885_ _06885_/A VGND VGND VPWR VPWR _07947_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _08645_/A _08505_/X _08546_/Y VGND VGND VPWR VPWR _08624_/X sky130_fd_sc_hd__o21ba_1
XFILLER_55_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _09407_/B _09407_/C VGND VGND VPWR VPWR _08556_/B sky130_fd_sc_hd__and2_1
XFILLER_70_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07506_ _09258_/B VGND VGND VPWR VPWR _09257_/B sky130_fd_sc_hd__buf_2
XFILLER_50_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08486_ _08464_/X _08481_/Y _08485_/X VGND VGND VPWR VPWR _13437_/D sky130_fd_sc_hd__a21o_1
XFILLER_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07437_ _07399_/X _07434_/Y _07436_/Y VGND VGND VPWR VPWR _13144_/D sky130_fd_sc_hd__a21o_1
XFILLER_22_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07368_ _07338_/X _07367_/Y _07355_/A VGND VGND VPWR VPWR _07369_/B sky130_fd_sc_hd__a21o_1
XFILLER_136_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09107_ _13527_/Q _09113_/B VGND VGND VPWR VPWR _09109_/B sky130_fd_sc_hd__xnor2_1
X_06319_ _14186_/D _14187_/D _06319_/C VGND VGND VPWR VPWR _06319_/Y sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_111_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _13606_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_108_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07299_ _13661_/Q _13659_/Q _07299_/S VGND VGND VPWR VPWR _07299_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09038_ _13219_/Q _13448_/Q _09040_/S VGND VGND VPWR VPWR _09039_/A sky130_fd_sc_hd__mux2_1
Xhold360 hold360/A VGND VGND VPWR VPWR hold360/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold371 hold371/A VGND VGND VPWR VPWR hold371/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_105_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold382 hold382/A VGND VGND VPWR VPWR hold382/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_11000_ _14600_/Q _14562_/Q _14493_/Q _14445_/Q _10969_/X _10970_/X VGND VGND VPWR
+ VPWR _11001_/A sky130_fd_sc_hd__mux4_1
Xhold393 hold393/A VGND VGND VPWR VPWR hold393/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12951_ _13574_/CLK _12951_/D VGND VGND VPWR VPWR hold284/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_178_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _14707_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_58_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11902_ _11902_/A VGND VGND VPWR VPWR _14258_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _12885_/CLK _12882_/D hold1/X VGND VGND VPWR VPWR _12882_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _14645_/CLK _14621_/D VGND VGND VPWR VPWR hold131/A sky130_fd_sc_hd__dfxtp_4
XFILLER_27_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11833_ _11833_/A VGND VGND VPWR VPWR _14108_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14552_ _14724_/CLK _14552_/D VGND VGND VPWR VPWR _14552_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _11370_/X _14073_/Q _11766_/S VGND VGND VPWR VPWR _11765_/A sky130_fd_sc_hd__mux2_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13503_ _13855_/CLK hold271/X VGND VGND VPWR VPWR _13503_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _10715_/A VGND VGND VPWR VPWR _12935_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14483_ _14510_/CLK _14483_/D VGND VGND VPWR VPWR _14483_/Q sky130_fd_sc_hd__dfxtp_1
X_11695_ _11695_/A VGND VGND VPWR VPWR _14029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13434_ _13434_/CLK hold210/X VGND VGND VPWR VPWR _13434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10646_ _14382_/Q _10646_/B VGND VGND VPWR VPWR _14358_/D sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_102_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _13686_/CLK sky130_fd_sc_hd__clkbuf_16
X_13365_ _13366_/CLK _13365_/D repeater56/X VGND VGND VPWR VPWR _13365_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10577_ _10510_/B _10521_/B _10576_/Y VGND VGND VPWR VPWR _14432_/D sky130_fd_sc_hd__a21oi_1
XFILLER_10_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12316_ _14573_/Q _12000_/X _12324_/S VGND VGND VPWR VPWR _12317_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13296_ _13296_/CLK hold19/X VGND VGND VPWR VPWR _13296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12247_ _12247_/A VGND VGND VPWR VPWR _14539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12178_ _12178_/A VGND VGND VPWR VPWR _14500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11129_ _14609_/Q _14571_/Q _14502_/Q _14454_/Q _11115_/X _11116_/X VGND VGND VPWR
+ VPWR _11130_/A sky130_fd_sc_hd__mux4_1
XFILLER_84_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_169_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _14424_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06670_ _06852_/B _06668_/X _06783_/S VGND VGND VPWR VPWR _06799_/B sky130_fd_sc_hd__mux2_1
XFILLER_36_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08340_ _13381_/Q _13384_/Q _08340_/C _08340_/D VGND VGND VPWR VPWR _08340_/X sky130_fd_sc_hd__and4_1
XFILLER_149_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08271_ _13368_/Q _08272_/B VGND VGND VPWR VPWR _08273_/A sky130_fd_sc_hd__and2_1
X_07222_ _07791_/A VGND VGND VPWR VPWR _13169_/D sky130_fd_sc_hd__clkbuf_2
X_07153_ _07153_/A _07153_/B _07153_/C VGND VGND VPWR VPWR _07155_/A sky130_fd_sc_hd__or3_1
XFILLER_146_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06104_ _06104_/A VGND VGND VPWR VPWR _13942_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07084_ hold187/A hold515/A _13708_/Q _14630_/Q VGND VGND VPWR VPWR _07114_/A sky130_fd_sc_hd__and4_1
XFILLER_160_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06035_ _06035_/A VGND VGND VPWR VPWR _06371_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_114_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07986_ _07986_/A _07986_/B VGND VGND VPWR VPWR _07987_/B sky130_fd_sc_hd__and2_1
XFILLER_68_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09725_ _09725_/A _09725_/B VGND VGND VPWR VPWR _09726_/B sky130_fd_sc_hd__or2_1
X_06937_ _06874_/X _06936_/Y _06897_/X VGND VGND VPWR VPWR _13019_/D sky130_fd_sc_hd__a21o_1
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09656_ _09656_/A VGND VGND VPWR VPWR _12840_/D sky130_fd_sc_hd__buf_2
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06868_ _06868_/A _06868_/B VGND VGND VPWR VPWR _06876_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08607_ _08607_/A _08607_/B _08607_/C VGND VGND VPWR VPWR _08671_/C sky130_fd_sc_hd__or3_1
XFILLER_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ _13392_/Q _13590_/Q _09587_/S VGND VGND VPWR VPWR _09588_/A sky130_fd_sc_hd__mux2_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06799_ _06863_/A _06799_/B VGND VGND VPWR VPWR _06800_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _13441_/Q _09399_/B VGND VGND VPWR VPWR _08538_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_23_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08469_ _08645_/B _08467_/X _08579_/S VGND VGND VPWR VPWR _08595_/B sky130_fd_sc_hd__mux2_1
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10500_ _10500_/A VGND VGND VPWR VPWR _14011_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11480_ _11480_/A VGND VGND VPWR VPWR _13828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10431_ _10431_/A _10431_/B VGND VGND VPWR VPWR _14440_/D sky130_fd_sc_hd__nand2_1
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13150_ _13555_/CLK _13150_/D repeater57/X VGND VGND VPWR VPWR _13150_/Q sky130_fd_sc_hd__dfrtp_1
X_10362_ _10386_/A VGND VGND VPWR VPWR _10415_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_151_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12101_ _12101_/A VGND VGND VPWR VPWR _14466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10293_ _10293_/A VGND VGND VPWR VPWR _12402_/B sky130_fd_sc_hd__clkbuf_1
X_13081_ _13434_/CLK hold121/X VGND VGND VPWR VPWR _13081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12032_ _14683_/Q _12034_/B VGND VGND VPWR VPWR _12033_/A sky130_fd_sc_hd__and2_1
XFILLER_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold190 hold190/A VGND VGND VPWR VPWR hold190/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13983_ _14705_/CLK _13983_/D VGND VGND VPWR VPWR _13983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12934_ _13265_/CLK _12934_/D VGND VGND VPWR VPWR hold369/A sky130_fd_sc_hd__dfxtp_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12865_ _13698_/CLK _12865_/D VGND VGND VPWR VPWR hold158/A sky130_fd_sc_hd__dfxtp_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _14605_/CLK _14604_/D VGND VGND VPWR VPWR _14604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _11816_/A VGND VGND VPWR VPWR _14100_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _13570_/CLK _12796_/D VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__dfxtp_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14535_ _14535_/CLK _14535_/D VGND VGND VPWR VPWR _14535_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11326_/X _14065_/Q _11747_/S VGND VGND VPWR VPWR _11748_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14466_ _14704_/CLK _14466_/D VGND VGND VPWR VPWR _14466_/Q sky130_fd_sc_hd__dfxtp_1
X_11678_ _14022_/Q _11478_/X _11678_/S VGND VGND VPWR VPWR _11679_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13417_ _14696_/CLK hold470/X VGND VGND VPWR VPWR _13417_/Q sky130_fd_sc_hd__dfxtp_1
X_10629_ _10206_/S _10626_/X _10627_/X _10628_/X _14383_/Q VGND VGND VPWR VPWR _14425_/D
+ sky130_fd_sc_hd__a221o_1
X_14397_ _14397_/CLK _14397_/D VGND VGND VPWR VPWR _14397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13348_ _14432_/CLK _13348_/D VGND VGND VPWR VPWR _13348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13279_ _13314_/CLK _13279_/D repeater59/X VGND VGND VPWR VPWR _13279_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07840_ _13257_/Q _07840_/B VGND VGND VPWR VPWR _07840_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07771_ _07772_/B _07785_/C _07785_/B _07772_/A VGND VGND VPWR VPWR _07773_/A sky130_fd_sc_hd__a22oi_1
XFILLER_77_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09510_ _09510_/A _09535_/A VGND VGND VPWR VPWR _09510_/X sky130_fd_sc_hd__or2_1
X_06722_ _06733_/B _06737_/A VGND VGND VPWR VPWR _06723_/A sky130_fd_sc_hd__and2_1
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09441_ _09448_/C _09448_/D VGND VGND VPWR VPWR _09454_/D sky130_fd_sc_hd__or2_1
X_06653_ _06690_/A VGND VGND VPWR VPWR _07804_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09372_ _08454_/X _09371_/X _09404_/S VGND VGND VPWR VPWR _09373_/A sky130_fd_sc_hd__mux2_1
X_06584_ _12894_/Q _12895_/Q _06584_/C _06584_/D VGND VGND VPWR VPWR _06598_/C sky130_fd_sc_hd__and4_1
XFILLER_33_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08323_ _13379_/Q _08322_/A _08298_/X VGND VGND VPWR VPWR _08323_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08254_ _08254_/A VGND VGND VPWR VPWR _08257_/A sky130_fd_sc_hd__inv_2
XFILLER_137_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07205_ _07205_/A _07205_/B _07205_/C VGND VGND VPWR VPWR _07206_/B sky130_fd_sc_hd__and3_1
X_08185_ _08261_/A _14012_/Q _08197_/A _08177_/A VGND VGND VPWR VPWR _08186_/C sky130_fd_sc_hd__a31o_1
XFILLER_119_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07136_ _07156_/A _07136_/B VGND VGND VPWR VPWR _07136_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_146_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07067_ _07067_/A _07067_/B VGND VGND VPWR VPWR _07069_/A sky130_fd_sc_hd__nor2_1
X_06018_ _13563_/Q _13574_/Q _06018_/C _06018_/D VGND VGND VPWR VPWR _06019_/B sky130_fd_sc_hd__or4_1
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07969_ _07970_/A _07970_/B _07970_/C VGND VGND VPWR VPWR _07969_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_101_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09708_ _09725_/A _09708_/B VGND VGND VPWR VPWR _09711_/A sky130_fd_sc_hd__or2_1
XFILLER_28_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10980_ _14298_/Q _14468_/Q _14224_/Q _14054_/Q _10914_/X _12643_/A VGND VGND VPWR
+ VPWR _10980_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09639_ _09639_/A VGND VGND VPWR VPWR _12832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12650_ _14744_/Q _12567_/X _12649_/X _12609_/X VGND VGND VPWR VPWR _14749_/D sky130_fd_sc_hd__o211a_1
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11601_ _12226_/A _12428_/B VGND VGND VPWR VPWR _11636_/A sky130_fd_sc_hd__nor2_8
X_12581_ _12619_/B _12578_/X _12580_/X VGND VGND VPWR VPWR _14727_/D sky130_fd_sc_hd__o21ai_1
X_14320_ _14357_/CLK hold114/X VGND VGND VPWR VPWR _14320_/Q sky130_fd_sc_hd__dfxtp_1
X_11532_ _11591_/B VGND VGND VPWR VPWR _11541_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_11_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14251_ _14251_/CLK _14251_/D VGND VGND VPWR VPWR _14251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11463_ _13823_/Q _11462_/X _11463_/S VGND VGND VPWR VPWR _11464_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13202_ _13372_/CLK _13202_/D VGND VGND VPWR VPWR hold66/A sky130_fd_sc_hd__dfxtp_1
X_10414_ _10415_/A _10429_/C _10415_/C VGND VGND VPWR VPWR _10416_/A sky130_fd_sc_hd__a21oi_1
XFILLER_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14182_ _14196_/CLK _14182_/D VGND VGND VPWR VPWR _14182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11394_ _13721_/Q _11394_/B VGND VGND VPWR VPWR _11395_/A sky130_fd_sc_hd__and2_1
XFILLER_99_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13133_ _13524_/CLK _13133_/D hold1/X VGND VGND VPWR VPWR _13133_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10345_ _10345_/A VGND VGND VPWR VPWR _13120_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_125_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _14082_/CLK _13064_/D VGND VGND VPWR VPWR hold139/A sky130_fd_sc_hd__dfxtp_1
X_10276_ _10286_/S VGND VGND VPWR VPWR _10592_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_155_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12015_ _12015_/A VGND VGND VPWR VPWR _14314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13966_ _13978_/CLK _13966_/D VGND VGND VPWR VPWR _13966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12917_ _14710_/CLK _12917_/D VGND VGND VPWR VPWR hold306/A sky130_fd_sc_hd__dfxtp_1
X_13897_ _14657_/CLK hold25/X VGND VGND VPWR VPWR hold371/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12848_ _13721_/CLK _12848_/D VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _13574_/CLK _12779_/D VGND VGND VPWR VPWR hold178/A sky130_fd_sc_hd__dfxtp_1
XFILLER_148_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14518_ _14716_/CLK _14518_/D VGND VGND VPWR VPWR _14518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14449_ _14712_/CLK _14449_/D VGND VGND VPWR VPWR _14449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09990_ _14428_/Q _14593_/Q _10597_/A VGND VGND VPWR VPWR _09990_/X sky130_fd_sc_hd__mux2_1
X_08941_ _08941_/A _08941_/B _08941_/C VGND VGND VPWR VPWR _08943_/A sky130_fd_sc_hd__or3_1
XFILLER_130_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08872_ _14003_/Q _13428_/Q _13519_/D _13520_/D VGND VGND VPWR VPWR _08902_/A sky130_fd_sc_hd__and4_1
XFILLER_69_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07823_ _07823_/A _07823_/B VGND VGND VPWR VPWR _07823_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_85_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07754_ _07721_/A _07785_/B _07729_/B _07753_/X VGND VGND VPWR VPWR _07756_/B sky130_fd_sc_hd__a31oi_1
X_06705_ _13348_/Q _13346_/Q _06705_/S VGND VGND VPWR VPWR _06705_/X sky130_fd_sc_hd__mux2_1
X_07685_ _07800_/S VGND VGND VPWR VPWR _07781_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_25_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_91_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _14251_/CLK sky130_fd_sc_hd__clkbuf_16
X_09424_ _13598_/Q _09424_/B _09424_/C VGND VGND VPWR VPWR _09447_/C sky130_fd_sc_hd__and3_1
X_06636_ _13034_/Q _13039_/Q VGND VGND VPWR VPWR _06636_/Y sky130_fd_sc_hd__nor2_2
XFILLER_12_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09355_ _09355_/A VGND VGND VPWR VPWR _12803_/D sky130_fd_sc_hd__clkbuf_1
X_06567_ _06567_/A VGND VGND VPWR VPWR _06567_/Y sky130_fd_sc_hd__inv_2
X_08306_ _08306_/A VGND VGND VPWR VPWR _13373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09286_ _09287_/B _09287_/C _09287_/A VGND VGND VPWR VPWR _09286_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06498_ _06499_/A _06499_/C _06499_/B VGND VGND VPWR VPWR _06498_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08237_ _08237_/A _08237_/B VGND VGND VPWR VPWR _08237_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_147_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08168_ _08137_/A _08136_/A _08152_/X _08151_/B VGND VGND VPWR VPWR _08169_/B sky130_fd_sc_hd__a211oi_1
XFILLER_109_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07119_ _07119_/A _07119_/B hold154/A _13115_/D VGND VGND VPWR VPWR _07150_/A sky130_fd_sc_hd__and4_1
X_08099_ _08099_/A VGND VGND VPWR VPWR _12708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10130_ _10130_/A VGND VGND VPWR VPWR _14179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10061_ _13918_/Q _10056_/X _10063_/A VGND VGND VPWR VPWR _14041_/D sky130_fd_sc_hd__a21o_1
XFILLER_88_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13820_ _14725_/CLK _13820_/D VGND VGND VPWR VPWR _13820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13751_ _14633_/CLK _13751_/D VGND VGND VPWR VPWR hold136/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10963_ _13319_/Q _10907_/X _10953_/X _10962_/Y VGND VGND VPWR VPWR _13319_/D sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_82_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _14687_/CLK sky130_fd_sc_hd__clkbuf_16
X_12702_ _14275_/CLK _12702_/D VGND VGND VPWR VPWR hold448/A sky130_fd_sc_hd__dfxtp_1
X_13682_ _13727_/CLK _13682_/D repeater56/X VGND VGND VPWR VPWR _13682_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10894_ _10894_/A VGND VGND VPWR VPWR _13205_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12633_ _12635_/B _12633_/B _12633_/C VGND VGND VPWR VPWR _12634_/A sky130_fd_sc_hd__and3b_1
XFILLER_43_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12564_ _12564_/A VGND VGND VPWR VPWR _12623_/B sky130_fd_sc_hd__clkbuf_2
X_14303_ _14495_/CLK _14303_/D VGND VGND VPWR VPWR _14303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11515_ _11515_/A VGND VGND VPWR VPWR _13839_/D sky130_fd_sc_hd__clkbuf_1
X_12495_ _12495_/A VGND VGND VPWR VPWR _14677_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14234_ _14652_/CLK _14234_/D VGND VGND VPWR VPWR _14234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11446_ _14694_/Q VGND VGND VPWR VPWR _11446_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14165_ _14209_/CLK hold390/X VGND VGND VPWR VPWR _14165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11377_ _11377_/A VGND VGND VPWR VPWR _13778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13116_ _13666_/CLK _13116_/D VGND VGND VPWR VPWR _13116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10328_ _13108_/Q _13241_/D VGND VGND VPWR VPWR _10329_/B sky130_fd_sc_hd__xor2_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _14397_/CLK _14096_/D VGND VGND VPWR VPWR _14096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _13528_/CLK _13047_/D VGND VGND VPWR VPWR hold138/A sky130_fd_sc_hd__dfxtp_1
X_10259_ _10190_/A _10237_/X _10246_/X VGND VGND VPWR VPWR _10259_/X sky130_fd_sc_hd__a21o_1
XFILLER_79_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13949_ _13964_/CLK _13949_/D VGND VGND VPWR VPWR _13949_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_73_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _13596_/CLK sky130_fd_sc_hd__clkbuf_16
X_07470_ _09270_/B VGND VGND VPWR VPWR _09277_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06421_ _06421_/A _06436_/A _06421_/C VGND VGND VPWR VPWR _06421_/X sky130_fd_sc_hd__and3_1
XFILLER_50_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09140_ _13532_/Q _09140_/B VGND VGND VPWR VPWR _09161_/C sky130_fd_sc_hd__nor2_1
X_06352_ _14403_/D _14404_/D _06348_/X _06351_/Y VGND VGND VPWR VPWR _14410_/D sky130_fd_sc_hd__a31o_1
XFILLER_148_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06283_ hold52/A _13952_/D _13954_/D _13955_/D VGND VGND VPWR VPWR _06284_/D sky130_fd_sc_hd__or4_1
X_09071_ _13233_/Q _13462_/Q _09075_/S VGND VGND VPWR VPWR _09072_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08022_ _08016_/A _08017_/X _08020_/Y _06859_/A VGND VGND VPWR VPWR _08022_/X sky130_fd_sc_hd__a31o_1
XFILLER_116_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09973_ _09973_/A VGND VGND VPWR VPWR _12872_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08924_ _08944_/A _08924_/B VGND VGND VPWR VPWR _08924_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_131_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08855_ _08855_/A _08855_/B VGND VGND VPWR VPWR _08857_/A sky130_fd_sc_hd__nor2_1
X_07806_ _07806_/A _07805_/X VGND VGND VPWR VPWR _07808_/A sky130_fd_sc_hd__or2b_1
XFILLER_57_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08786_ _08786_/A _08786_/B _08779_/Y _08780_/X VGND VGND VPWR VPWR _08791_/C sky130_fd_sc_hd__or4bb_1
X_05998_ _10224_/S VGND VGND VPWR VPWR _14384_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07737_ _07737_/A _07764_/B VGND VGND VPWR VPWR _07738_/B sky130_fd_sc_hd__nand2_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_64_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _13528_/CLK sky130_fd_sc_hd__clkbuf_16
X_07668_ _07665_/Y _07696_/A _07668_/C _13246_/D VGND VGND VPWR VPWR _07696_/B sky130_fd_sc_hd__and4bb_1
XFILLER_53_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09407_ _13596_/Q _09407_/B _09407_/C VGND VGND VPWR VPWR _09420_/A sky130_fd_sc_hd__and3_1
X_06619_ _12904_/Q _12905_/Q _12906_/Q VGND VGND VPWR VPWR _06620_/C sky130_fd_sc_hd__and3_1
XFILLER_25_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07599_ _13244_/D _07645_/B VGND VGND VPWR VPWR _07627_/C sky130_fd_sc_hd__and2_1
XFILLER_13_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09338_ _09338_/A VGND VGND VPWR VPWR _12795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09269_ _09256_/A _09256_/B _09267_/Y _09268_/X VGND VGND VPWR VPWR _09282_/A sky130_fd_sc_hd__a31oi_2
X_11300_ _11300_/A VGND VGND VPWR VPWR _13760_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12280_ _12428_/B _12342_/B VGND VGND VPWR VPWR _12315_/A sky130_fd_sc_hd__nor2_4
XFILLER_4_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11231_ _11242_/A _11231_/B VGND VGND VPWR VPWR _11231_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11162_ _11162_/A VGND VGND VPWR VPWR _11162_/X sky130_fd_sc_hd__buf_2
XFILLER_150_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10113_ _10616_/C _10111_/X _10119_/S VGND VGND VPWR VPWR _10114_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11093_ _14267_/Q _14658_/Q _13765_/Q _14713_/Q _11091_/X _11092_/X VGND VGND VPWR
+ VPWR _11094_/B sky130_fd_sc_hd__mux4_1
XFILLER_122_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10044_ _13802_/Q _13786_/Q _13935_/D VGND VGND VPWR VPWR _10045_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_102_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold61 hold61/A VGND VGND VPWR VPWR hold61/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold72 hold72/A VGND VGND VPWR VPWR hold72/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold83 hold83/A VGND VGND VPWR VPWR hold83/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold94 hold94/A VGND VGND VPWR VPWR hold94/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_91_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13803_ _13843_/CLK _13803_/D VGND VGND VPWR VPWR _13803_/Q sky130_fd_sc_hd__dfxtp_1
X_11995_ _14308_/Q _11994_/X _11998_/S VGND VGND VPWR VPWR _11996_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _14644_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13734_ _13805_/CLK hold231/X VGND VGND VPWR VPWR _13734_/Q sky130_fd_sc_hd__dfxtp_1
X_10946_ _11224_/A VGND VGND VPWR VPWR _10946_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13665_ _13666_/CLK _13665_/D VGND VGND VPWR VPWR _13665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10877_ _13155_/Q _10885_/B VGND VGND VPWR VPWR _10878_/A sky130_fd_sc_hd__and2_1
XFILLER_31_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12616_ _12616_/A _12616_/B VGND VGND VPWR VPWR _12616_/X sky130_fd_sc_hd__or2_1
X_13596_ _13596_/CLK _13596_/D repeater56/X VGND VGND VPWR VPWR _13596_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12547_ _12547_/A VGND VGND VPWR VPWR _14718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12478_ _14670_/Q _12022_/A _12480_/S VGND VGND VPWR VPWR _12479_/A sky130_fd_sc_hd__mux2_1
XANTENNA_3 _11636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14217_ _14440_/CLK _14217_/D VGND VGND VPWR VPWR _14217_/Q sky130_fd_sc_hd__dfxtp_1
X_11429_ _11429_/A VGND VGND VPWR VPWR _11438_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14148_ _14153_/CLK _14148_/D VGND VGND VPWR VPWR hold184/A sky130_fd_sc_hd__dfxtp_1
XFILLER_141_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14079_ _14397_/CLK _14079_/D VGND VGND VPWR VPWR _14079_/Q sky130_fd_sc_hd__dfxtp_1
X_06970_ _13024_/Q _07989_/B VGND VGND VPWR VPWR _06971_/B sky130_fd_sc_hd__or2_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05921_ _13843_/D _13721_/Q _05921_/C _05921_/D VGND VGND VPWR VPWR _05921_/Y sky130_fd_sc_hd__nor4_1
XFILLER_66_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08640_ _13447_/Q _09450_/B _08629_/X VGND VGND VPWR VPWR _08644_/B sky130_fd_sc_hd__a21bo_1
XFILLER_54_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08571_ _13443_/Q _08577_/B VGND VGND VPWR VPWR _08622_/A sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_46_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _14692_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_82_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07522_ _07530_/A _07522_/B VGND VGND VPWR VPWR _07532_/C sky130_fd_sc_hd__or2_1
XFILLER_23_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07453_ _07454_/A _07454_/B _07454_/C VGND VGND VPWR VPWR _07453_/X sky130_fd_sc_hd__a21o_1
XFILLER_62_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06404_ _06471_/A VGND VGND VPWR VPWR _10349_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_07384_ _09140_/B _07383_/Y _09182_/A VGND VGND VPWR VPWR _07385_/A sky130_fd_sc_hd__mux2_1
X_09123_ _09134_/C _09122_/B _07341_/A VGND VGND VPWR VPWR _09123_/Y sky130_fd_sc_hd__a21oi_1
X_06335_ _14104_/Q _14088_/Q _06345_/S VGND VGND VPWR VPWR _06336_/A sky130_fd_sc_hd__mux2_1
X_09054_ _09644_/A VGND VGND VPWR VPWR _09600_/A sky130_fd_sc_hd__buf_2
X_06266_ _13806_/Q _13790_/Q _06273_/S VGND VGND VPWR VPWR _06267_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08005_ _08013_/A _08013_/B _06836_/X VGND VGND VPWR VPWR _08005_/X sky130_fd_sc_hd__a21o_1
Xhold520 hold520/A VGND VGND VPWR VPWR hold520/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_06197_ _06197_/A VGND VGND VPWR VPWR _10193_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09956_ _09956_/A VGND VGND VPWR VPWR _12864_/D sky130_fd_sc_hd__clkbuf_1
X_08907_ _08907_/A _08907_/B _13431_/Q _13432_/Q VGND VGND VPWR VPWR _08938_/A sky130_fd_sc_hd__and4_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _13694_/Q _09885_/B _09855_/X VGND VGND VPWR VPWR _09888_/B sky130_fd_sc_hd__o21ai_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08838_ _08816_/B _08820_/B _08816_/A VGND VGND VPWR VPWR _08839_/B sky130_fd_sc_hd__o21ba_1
XFILLER_100_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ _08633_/X _08768_/Y _08684_/X VGND VGND VPWR VPWR _13462_/D sky130_fd_sc_hd__a21o_1
XFILLER_72_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _12930_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _10800_/A VGND VGND VPWR VPWR _13062_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _13562_/Q _11784_/B VGND VGND VPWR VPWR _11781_/A sky130_fd_sc_hd__and2_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10731_ _12900_/Q _10731_/B VGND VGND VPWR VPWR _10732_/A sky130_fd_sc_hd__and2_1
XFILLER_14_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13450_ _13602_/CLK _13450_/D repeater57/X VGND VGND VPWR VPWR _13450_/Q sky130_fd_sc_hd__dfrtp_1
X_10662_ _10662_/A VGND VGND VPWR VPWR _12913_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12401_ _12401_/A VGND VGND VPWR VPWR hold461/A sky130_fd_sc_hd__clkbuf_1
X_13381_ _14333_/CLK _13381_/D _12609_/A VGND VGND VPWR VPWR _13381_/Q sky130_fd_sc_hd__dfrtp_1
X_10593_ _10593_/A _14583_/Q VGND VGND VPWR VPWR _13747_/D sky130_fd_sc_hd__xor2_1
X_12332_ _14581_/Q _12025_/X _12332_/S VGND VGND VPWR VPWR _12333_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12263_ _12263_/A VGND VGND VPWR VPWR _14546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14002_ _14725_/CLK _14002_/D VGND VGND VPWR VPWR _14002_/Q sky130_fd_sc_hd__dfxtp_1
X_11214_ _14615_/Q _14577_/Q _14508_/Q _14460_/Q _11186_/X _11187_/X VGND VGND VPWR
+ VPWR _11215_/A sky130_fd_sc_hd__mux4_1
X_12194_ _14508_/Q _12013_/X _12194_/S VGND VGND VPWR VPWR _12195_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput40 _13337_/Q VGND VGND VPWR VPWR data_o[19] sky130_fd_sc_hd__buf_2
Xoutput51 _13325_/Q VGND VGND VPWR VPWR data_o[7] sky130_fd_sc_hd__buf_2
XFILLER_150_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11145_ _14271_/Q _14662_/Q _13769_/Q _14717_/Q _11091_/X _11092_/X VGND VGND VPWR
+ VPWR _11146_/B sky130_fd_sc_hd__mux4_1
XFILLER_150_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11076_ _11017_/X _11073_/Y _11075_/Y _11024_/X VGND VGND VPWR VPWR _11077_/B sky130_fd_sc_hd__a211o_1
XFILLER_48_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10027_ _10027_/A VGND VGND VPWR VPWR _13968_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_28_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _13296_/CLK sky130_fd_sc_hd__clkbuf_16
X_11978_ _14513_/Q VGND VGND VPWR VPWR _11978_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10929_ _10929_/A VGND VGND VPWR VPWR _10929_/X sky130_fd_sc_hd__clkbuf_2
X_13717_ _13799_/CLK hold137/X VGND VGND VPWR VPWR _13717_/Q sky130_fd_sc_hd__dfxtp_1
X_14697_ _14697_/CLK hold238/X VGND VGND VPWR VPWR _14697_/Q sky130_fd_sc_hd__dfxtp_2
X_13648_ _14327_/CLK hold396/X VGND VGND VPWR VPWR _13648_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13579_ _14319_/CLK hold50/X VGND VGND VPWR VPWR _13579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06120_ _06116_/X _06117_/X _06127_/A VGND VGND VPWR VPWR _06121_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06051_ _06051_/A VGND VGND VPWR VPWR _13916_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09810_ _13679_/Q _09811_/B VGND VGND VPWR VPWR _09812_/A sky130_fd_sc_hd__and2_1
XFILLER_113_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09741_ _09741_/A _09741_/B VGND VGND VPWR VPWR _09741_/X sky130_fd_sc_hd__xor2_1
XFILLER_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06953_ _06899_/A _06951_/Y _06952_/X _06926_/X VGND VGND VPWR VPWR _06968_/A sky130_fd_sc_hd__a211o_2
XFILLER_28_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05904_ _13800_/Q _13801_/Q _05904_/C _05904_/D VGND VGND VPWR VPWR _05911_/A sky130_fd_sc_hd__nor4_1
X_09672_ _13701_/Q VGND VGND VPWR VPWR _09672_/Y sky130_fd_sc_hd__inv_2
X_06884_ _13014_/Q _07955_/B VGND VGND VPWR VPWR _06887_/A sky130_fd_sc_hd__nand2_1
XFILLER_94_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08623_ _08539_/X _08572_/Y _08621_/C _08622_/X _08558_/A VGND VGND VPWR VPWR _08630_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_54_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _13587_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08554_ _08567_/A _08552_/A _08552_/B _08552_/C VGND VGND VPWR VPWR _09407_/C sky130_fd_sc_hd__a31o_1
XFILLER_35_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07505_ _07533_/A VGND VGND VPWR VPWR _07505_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08485_ _08642_/A _09383_/B VGND VGND VPWR VPWR _08485_/X sky130_fd_sc_hd__and2_1
XFILLER_23_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07436_ _09125_/A _09177_/B VGND VGND VPWR VPWR _07436_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07367_ _07367_/A _07367_/B VGND VGND VPWR VPWR _07367_/Y sky130_fd_sc_hd__nor2_1
X_09106_ _09182_/A VGND VGND VPWR VPWR _09106_/X sky130_fd_sc_hd__clkbuf_2
X_06318_ _14189_/D _14190_/D _14191_/D _06318_/D VGND VGND VPWR VPWR _06319_/C sky130_fd_sc_hd__or4_1
XFILLER_148_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07298_ _13665_/Q _13663_/Q _07299_/S VGND VGND VPWR VPWR _07298_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09037_ _09037_/A VGND VGND VPWR VPWR _12754_/D sky130_fd_sc_hd__clkbuf_1
X_06249_ _14083_/Q _14084_/Q _14085_/Q _14086_/Q VGND VGND VPWR VPWR _06249_/X sky130_fd_sc_hd__or4_1
XFILLER_105_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold350 hold350/A VGND VGND VPWR VPWR hold350/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold361 hold361/A VGND VGND VPWR VPWR hold361/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold372 hold372/A VGND VGND VPWR VPWR hold372/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold383 hold383/A VGND VGND VPWR VPWR hold383/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold394 hold394/A VGND VGND VPWR VPWR hold394/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_120_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09939_ _09939_/A VGND VGND VPWR VPWR _12856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_13_0_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR clkbuf_4_13_0_clk/X sky130_fd_sc_hd__clkbuf_2
X_12950_ _13274_/CLK _12950_/D VGND VGND VPWR VPWR hold333/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11901_ _14258_/Q _11453_/X _11907_/S VGND VGND VPWR VPWR _11902_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _12881_/CLK _12881_/D hold1/X VGND VGND VPWR VPWR _12881_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _13586_/Q _11834_/B VGND VGND VPWR VPWR _11833_/A sky130_fd_sc_hd__and2_1
XFILLER_73_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14620_ _14679_/CLK _14646_/Q VGND VGND VPWR VPWR hold205/A sky130_fd_sc_hd__dfxtp_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _14724_/CLK _14551_/D VGND VGND VPWR VPWR _14551_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _11763_/A VGND VGND VPWR VPWR _14072_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13502_ _13698_/CLK hold262/X VGND VGND VPWR VPWR _13502_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _12892_/Q _10720_/B VGND VGND VPWR VPWR _10715_/A sky130_fd_sc_hd__and2_1
X_14482_ _14510_/CLK _14482_/D VGND VGND VPWR VPWR _14482_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _14029_/Q _11501_/X _11700_/S VGND VGND VPWR VPWR _11695_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13433_ _14588_/CLK hold212/X VGND VGND VPWR VPWR _13433_/Q sky130_fd_sc_hd__dfxtp_1
X_10645_ _14411_/Q hold354/A _14385_/Q VGND VGND VPWR VPWR _10646_/B sky130_fd_sc_hd__o21ai_1
XFILLER_9_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13364_ _13366_/CLK _13364_/D repeater56/X VGND VGND VPWR VPWR _13364_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10576_ _10510_/B _10521_/B _10512_/A VGND VGND VPWR VPWR _10576_/Y sky130_fd_sc_hd__o21ai_1
X_12315_ _12315_/A VGND VGND VPWR VPWR _12324_/S sky130_fd_sc_hd__buf_2
XFILLER_5_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13295_ _13298_/CLK hold240/X VGND VGND VPWR VPWR _13295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12246_ _11307_/X _14539_/Q _12248_/S VGND VGND VPWR VPWR _12247_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12177_ _14500_/Q _11988_/X _12183_/S VGND VGND VPWR VPWR _12178_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11128_ _11065_/X _11125_/X _11127_/X _11086_/X VGND VGND VPWR VPWR _11128_/X sky130_fd_sc_hd__o211a_1
X_11059_ _11059_/A VGND VGND VPWR VPWR _11059_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14749_ _14749_/CLK _14749_/D VGND VGND VPWR VPWR _14749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08270_ _10304_/A _08270_/B _08279_/D VGND VGND VPWR VPWR _08272_/B sky130_fd_sc_hd__and3_1
XFILLER_20_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07221_ _07796_/A VGND VGND VPWR VPWR _07791_/A sky130_fd_sc_hd__clkbuf_2
X_07152_ _07152_/A _07152_/B VGND VGND VPWR VPWR _07153_/C sky130_fd_sc_hd__xnor2_2
XFILLER_145_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06103_ _13796_/Q _06105_/B VGND VGND VPWR VPWR _06104_/A sky130_fd_sc_hd__and2_1
XFILLER_145_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07083_ hold515/A _13708_/Q _14630_/Q _07063_/A VGND VGND VPWR VPWR _07083_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _13280_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_160_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06034_ input28/X input29/X VGND VGND VPWR VPWR _06035_/A sky130_fd_sc_hd__and2_1
XFILLER_160_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07985_ _13276_/Q _13277_/Q _06895_/B VGND VGND VPWR VPWR _07992_/B sky130_fd_sc_hd__o21ai_1
XFILLER_86_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09724_ _09697_/A _09696_/A _09709_/X _09708_/B VGND VGND VPWR VPWR _09725_/B sky130_fd_sc_hd__a211oi_1
X_06936_ _06936_/A _06951_/C VGND VGND VPWR VPWR _06936_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_55_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09655_ _13423_/Q _13621_/Q _09655_/S VGND VGND VPWR VPWR _09656_/A sky130_fd_sc_hd__mux2_1
X_06867_ _13013_/Q _07911_/B VGND VGND VPWR VPWR _06868_/B sky130_fd_sc_hd__or2_1
XFILLER_103_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08606_ _08657_/A _08606_/B VGND VGND VPWR VPWR _08607_/C sky130_fd_sc_hd__nor2_2
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_2_0_clk clkbuf_3_3_0_clk/A VGND VGND VPWR VPWR clkbuf_4_5_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_09586_ _09586_/A VGND VGND VPWR VPWR _12808_/D sky130_fd_sc_hd__clkbuf_2
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06798_ _06745_/X _06881_/B _06881_/A VGND VGND VPWR VPWR _06800_/A sky130_fd_sc_hd__o21ai_2
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _09399_/B VGND VGND VPWR VPWR _09417_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_11_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08468_ _13475_/Q VGND VGND VPWR VPWR _08579_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07419_ _07401_/A _07389_/B _07401_/C _07363_/B VGND VGND VPWR VPWR _07420_/A sky130_fd_sc_hd__o31a_1
XFILLER_156_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08399_ _08399_/A VGND VGND VPWR VPWR _12731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10430_ _10430_/A VGND VGND VPWR VPWR _14220_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10361_ _13517_/Q VGND VGND VPWR VPWR _10386_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12100_ _14466_/Q _11956_/X _12106_/S VGND VGND VPWR VPWR _12101_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13080_ _13434_/CLK hold138/X VGND VGND VPWR VPWR _13080_/Q sky130_fd_sc_hd__dfxtp_1
X_10292_ _13522_/Q VGND VGND VPWR VPWR _13701_/D sky130_fd_sc_hd__clkinv_2
XFILLER_105_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12031_ _12031_/A VGND VGND VPWR VPWR _14324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold180 hold180/A VGND VGND VPWR VPWR hold180/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold191 hold191/A VGND VGND VPWR VPWR hold191/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13982_ _14533_/CLK _13982_/D VGND VGND VPWR VPWR _13982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12933_ _13265_/CLK _12933_/D VGND VGND VPWR VPWR hold196/A sky130_fd_sc_hd__dfxtp_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12864_ _13700_/CLK _12864_/D VGND VGND VPWR VPWR hold130/A sky130_fd_sc_hd__dfxtp_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _14605_/CLK _14603_/D VGND VGND VPWR VPWR _14603_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _13578_/Q _11817_/B VGND VGND VPWR VPWR _11816_/A sky130_fd_sc_hd__and2_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _13570_/CLK _12795_/D VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__dfxtp_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _11746_/A VGND VGND VPWR VPWR _14064_/D sky130_fd_sc_hd__clkbuf_1
X_14534_ _14535_/CLK _14534_/D VGND VGND VPWR VPWR _14534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14465_ _14742_/CLK _14465_/D VGND VGND VPWR VPWR _14465_/Q sky130_fd_sc_hd__dfxtp_1
X_11677_ _11677_/A VGND VGND VPWR VPWR _14021_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10628_ _14413_/Q _14386_/Q _10627_/A VGND VGND VPWR VPWR _10628_/X sky130_fd_sc_hd__or3b_1
X_13416_ _14696_/CLK hold363/X VGND VGND VPWR VPWR _13416_/Q sky130_fd_sc_hd__dfxtp_1
X_14396_ _14413_/CLK _14396_/D VGND VGND VPWR VPWR _14396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13347_ _14680_/CLK _13347_/D VGND VGND VPWR VPWR _13347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10559_ _10557_/A _10573_/C _10526_/C _10547_/A _10545_/A VGND VGND VPWR VPWR _10560_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13278_ _13280_/CLK _13278_/D repeater59/X VGND VGND VPWR VPWR _13278_/Q sky130_fd_sc_hd__dfrtp_1
X_12229_ _11272_/X _14531_/Q _12237_/S VGND VGND VPWR VPWR _12230_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07770_ _07747_/A _07785_/B _07748_/A _07746_/B VGND VGND VPWR VPWR _07786_/A sky130_fd_sc_hd__a31o_1
XFILLER_84_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06721_ _06770_/A _06753_/A VGND VGND VPWR VPWR _06737_/A sky130_fd_sc_hd__nand2_2
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09440_ _13600_/Q _09440_/B _09440_/C VGND VGND VPWR VPWR _09448_/D sky130_fd_sc_hd__and3_1
X_06652_ _06736_/A _06881_/B _06652_/C _06652_/D VGND VGND VPWR VPWR _06690_/A sky130_fd_sc_hd__nand4_4
XFILLER_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09371_ _09371_/A _09371_/B VGND VGND VPWR VPWR _09371_/X sky130_fd_sc_hd__xor2_1
X_06583_ _06583_/A VGND VGND VPWR VPWR _12894_/D sky130_fd_sc_hd__clkbuf_1
X_08322_ _08322_/A _08322_/B VGND VGND VPWR VPWR _13378_/D sky130_fd_sc_hd__nor2_1
XFILLER_21_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08253_ _08253_/A _08253_/B VGND VGND VPWR VPWR _08254_/A sky130_fd_sc_hd__or2_1
XFILLER_119_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07204_ _07204_/A _07204_/B VGND VGND VPWR VPWR _07206_/A sky130_fd_sc_hd__and2_1
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08184_ _08114_/X _08126_/X _08129_/X _08162_/Y VGND VGND VPWR VPWR _08186_/B sky130_fd_sc_hd__o22a_1
XFILLER_20_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07135_ _07153_/B _07135_/B VGND VGND VPWR VPWR _07136_/B sky130_fd_sc_hd__or2_1
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07066_ hold425/A _13706_/Q _07086_/C hold177/A VGND VGND VPWR VPWR _07067_/B sky130_fd_sc_hd__and4_1
XFILLER_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06017_ _13572_/Q _13573_/Q _06017_/C _06017_/D VGND VGND VPWR VPWR _06018_/D sky130_fd_sc_hd__or4_1
XFILLER_133_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07968_ _13275_/Q _07968_/B VGND VGND VPWR VPWR _07970_/C sky130_fd_sc_hd__xor2_1
XFILLER_101_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06919_ _06919_/A _06919_/B _06924_/D VGND VGND VPWR VPWR _06919_/Y sky130_fd_sc_hd__nand3_1
X_09707_ _13670_/Q _09707_/B VGND VGND VPWR VPWR _09708_/B sky130_fd_sc_hd__and2_1
X_07899_ _07917_/A _07904_/B VGND VGND VPWR VPWR _07899_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09638_ _13415_/Q _13613_/Q _09642_/S VGND VGND VPWR VPWR _09639_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09569_ _13618_/Q _09569_/B VGND VGND VPWR VPWR _09569_/X sky130_fd_sc_hd__or2_1
X_11600_ _11655_/A _12614_/A _12582_/A VGND VGND VPWR VPWR _12428_/B sky130_fd_sc_hd__or3_4
X_12580_ _12641_/A VGND VGND VPWR VPWR _12580_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11531_ _11576_/A VGND VGND VPWR VPWR _11591_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_23_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14250_ _14250_/CLK _14250_/D VGND VGND VPWR VPWR _14250_/Q sky130_fd_sc_hd__dfxtp_1
X_11462_ _14698_/Q VGND VGND VPWR VPWR _11462_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13201_ _13617_/CLK _13201_/D VGND VGND VPWR VPWR hold426/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10413_ _10423_/A _10413_/B VGND VGND VPWR VPWR _10415_/C sky130_fd_sc_hd__and2_1
X_14181_ _14196_/CLK _14181_/D VGND VGND VPWR VPWR _14181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11393_ _11393_/A VGND VGND VPWR VPWR _13789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13132_ _13524_/CLK _13132_/D hold1/X VGND VGND VPWR VPWR _13132_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10344_ _10348_/B _10344_/B VGND VGND VPWR VPWR _10345_/A sky130_fd_sc_hd__or2_1
XFILLER_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ _13587_/CLK _13063_/D VGND VGND VPWR VPWR hold410/A sky130_fd_sc_hd__dfxtp_1
X_10275_ _14589_/Q _10275_/B VGND VGND VPWR VPWR _10286_/S sky130_fd_sc_hd__xnor2_1
XFILLER_124_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12014_ _14314_/Q _12013_/X _12014_/S VGND VGND VPWR VPWR _12015_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13965_ _14179_/CLK _13965_/D VGND VGND VPWR VPWR _13965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12916_ _14697_/CLK _12916_/D VGND VGND VPWR VPWR hold102/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13896_ _14050_/CLK hold148/X VGND VGND VPWR VPWR hold481/A sky130_fd_sc_hd__dfxtp_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _13727_/CLK _12847_/D VGND VGND VPWR VPWR hold179/A sky130_fd_sc_hd__dfxtp_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _13565_/CLK _12778_/D VGND VGND VPWR VPWR hold462/A sky130_fd_sc_hd__dfxtp_1
XFILLER_159_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14517_ _14608_/CLK _14517_/D VGND VGND VPWR VPWR _14517_/Q sky130_fd_sc_hd__dfxtp_1
X_11729_ _11729_/A VGND VGND VPWR VPWR _14056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14448_ _14712_/CLK _14448_/D VGND VGND VPWR VPWR _14448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14379_ _14732_/CLK hold77/X VGND VGND VPWR VPWR _14379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08940_ _08940_/A _08940_/B VGND VGND VPWR VPWR _08941_/C sky130_fd_sc_hd__xnor2_1
X_08871_ _13428_/Q _13519_/D _13520_/D _08851_/A VGND VGND VPWR VPWR _08871_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_130_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07822_ _07815_/A _07815_/B _07821_/X VGND VGND VPWR VPWR _07823_/B sky130_fd_sc_hd__a21o_1
XFILLER_85_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07753_ _07728_/B _07753_/B VGND VGND VPWR VPWR _07753_/X sky130_fd_sc_hd__and2b_1
XFILLER_37_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06704_ _13352_/Q _13350_/Q _06704_/S VGND VGND VPWR VPWR _06704_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07684_ _07738_/A _07684_/B VGND VGND VPWR VPWR _07684_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_38_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09423_ _09423_/A VGND VGND VPWR VPWR _13597_/D sky130_fd_sc_hd__clkbuf_1
X_06635_ _13352_/Q _13350_/Q _13348_/Q _13346_/Q _06704_/S _13038_/Q VGND VGND VPWR
+ VPWR _06767_/B sky130_fd_sc_hd__mux4_2
X_09354_ _13313_/Q _13551_/Q _09354_/S VGND VGND VPWR VPWR _09355_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06566_ _06566_/A _06566_/B VGND VGND VPWR VPWR _06569_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08305_ _08314_/B _09084_/A _08305_/C VGND VGND VPWR VPWR _08306_/A sky130_fd_sc_hd__and3b_1
X_09285_ _09285_/A _09285_/B VGND VGND VPWR VPWR _09287_/A sky130_fd_sc_hd__nand2_1
X_06497_ _12884_/Q _06500_/B VGND VGND VPWR VPWR _06499_/B sky130_fd_sc_hd__xnor2_1
XFILLER_20_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08236_ _08236_/A _08236_/B VGND VGND VPWR VPWR _08237_/B sky130_fd_sc_hd__and2_1
XFILLER_138_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08167_ _08167_/A _08167_/B VGND VGND VPWR VPWR _08170_/A sky130_fd_sc_hd__nand2_1
XFILLER_109_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07118_ _07139_/A _07190_/B _07190_/D _07119_/A VGND VGND VPWR VPWR _07120_/A sky130_fd_sc_hd__a22oi_1
XFILLER_106_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08098_ _12984_/Q _13284_/Q _10781_/A VGND VGND VPWR VPWR _08099_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07049_ _07059_/A _07049_/B VGND VGND VPWR VPWR _07058_/B sky130_fd_sc_hd__xnor2_1
XFILLER_122_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10060_ _10060_/A VGND VGND VPWR VPWR _10063_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13750_ _14432_/CLK _13750_/D VGND VGND VPWR VPWR _14430_/D sky130_fd_sc_hd__dfxtp_1
X_10962_ _10962_/A _10962_/B VGND VGND VPWR VPWR _10962_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12701_ _14275_/CLK _12701_/D VGND VGND VPWR VPWR hold368/A sky130_fd_sc_hd__dfxtp_1
X_10893_ _10893_/A _13163_/Q VGND VGND VPWR VPWR _10894_/A sky130_fd_sc_hd__and2_1
X_13681_ _13681_/CLK _13681_/D repeater56/X VGND VGND VPWR VPWR _13681_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_71_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12632_ _12631_/B _14740_/Q _11185_/A _14742_/Q VGND VGND VPWR VPWR _12633_/C sky130_fd_sc_hd__a31o_1
XFILLER_70_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12563_ _12563_/A VGND VGND VPWR VPWR _14726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14302_ _14495_/CLK _14302_/D VGND VGND VPWR VPWR _14302_/Q sky130_fd_sc_hd__dfxtp_1
X_11514_ _13839_/Q _11513_/X _11523_/S VGND VGND VPWR VPWR _11515_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12494_ _12496_/A _12496_/B hold150/X VGND VGND VPWR VPWR _12495_/A sky130_fd_sc_hd__and3_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14233_ _14543_/CLK _14233_/D VGND VGND VPWR VPWR _14233_/Q sky130_fd_sc_hd__dfxtp_1
X_11445_ _11445_/A VGND VGND VPWR VPWR _13813_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14164_ _14209_/CLK hold419/X VGND VGND VPWR VPWR hold390/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11376_ _13778_/Q _11375_/X _11376_/S VGND VGND VPWR VPWR _11377_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13115_ _14645_/CLK _13115_/D VGND VGND VPWR VPWR _13115_/Q sky130_fd_sc_hd__dfxtp_1
X_10327_ _10327_/A VGND VGND VPWR VPWR _13241_/D sky130_fd_sc_hd__buf_2
X_14095_ _14397_/CLK _14095_/D VGND VGND VPWR VPWR _14095_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _13528_/CLK _13046_/D VGND VGND VPWR VPWR hold122/A sky130_fd_sc_hd__dfxtp_1
X_10258_ _10258_/A VGND VGND VPWR VPWR _14352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10189_ _10226_/A _14361_/Q VGND VGND VPWR VPWR _10190_/A sky130_fd_sc_hd__xnor2_2
XFILLER_67_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13948_ _13964_/CLK _13948_/D VGND VGND VPWR VPWR _13948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13879_ _14657_/CLK hold334/X VGND VGND VPWR VPWR hold232/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06420_ _12878_/Q _06423_/B VGND VGND VPWR VPWR _06421_/C sky130_fd_sc_hd__nand2_1
X_06351_ _14403_/D _14404_/D _06351_/C VGND VGND VPWR VPWR _06351_/Y sky130_fd_sc_hd__nor3_1
X_09070_ _09070_/A VGND VGND VPWR VPWR _12768_/D sky130_fd_sc_hd__clkbuf_1
X_06282_ _06282_/A VGND VGND VPWR VPWR _13959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08021_ _08016_/A _08017_/X _08020_/Y VGND VGND VPWR VPWR _08021_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09972_ _13509_/Q _13698_/Q _09974_/S VGND VGND VPWR VPWR _09973_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08923_ _08941_/B _08923_/B VGND VGND VPWR VPWR _08924_/B sky130_fd_sc_hd__or2_1
XFILLER_69_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08854_ _13516_/D _13517_/D _08874_/C _13430_/Q VGND VGND VPWR VPWR _08855_/B sky130_fd_sc_hd__and4_1
XFILLER_84_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07805_ _07804_/B _07804_/C _13253_/Q VGND VGND VPWR VPWR _07805_/X sky130_fd_sc_hd__a21o_1
X_08785_ _13463_/Q _13464_/Q _09581_/B VGND VGND VPWR VPWR _08791_/B sky130_fd_sc_hd__o21ai_1
XFILLER_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05997_ _06345_/S VGND VGND VPWR VPWR _10224_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_85_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07736_ _07735_/A _07735_/B _07735_/C VGND VGND VPWR VPWR _07764_/B sky130_fd_sc_hd__o21ai_2
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07667_ _07668_/C _13246_/D _07665_/Y _07696_/A VGND VGND VPWR VPWR _07669_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_53_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06618_ _12905_/Q _06616_/A _06617_/Y VGND VGND VPWR VPWR _12905_/D sky130_fd_sc_hd__a21oi_1
XFILLER_80_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09406_ _09407_/B _09407_/C _13596_/Q VGND VGND VPWR VPWR _09408_/A sky130_fd_sc_hd__a21oi_1
XFILLER_25_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07598_ _07622_/A _07701_/A _07645_/B _07613_/A VGND VGND VPWR VPWR _07601_/A sky130_fd_sc_hd__a22oi_1
XFILLER_40_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09337_ _13305_/Q _13543_/Q _09343_/S VGND VGND VPWR VPWR _09338_/A sky130_fd_sc_hd__mux2_1
X_06549_ _06537_/A _06548_/Y _06537_/B _06535_/A VGND VGND VPWR VPWR _06550_/B sky130_fd_sc_hd__a31o_1
XFILLER_40_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09268_ _13547_/Q _13548_/Q _13549_/Q _13550_/Q _09271_/B VGND VGND VPWR VPWR _09268_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_138_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08219_ _13363_/Q _08220_/C _08250_/C VGND VGND VPWR VPWR _08222_/A sky130_fd_sc_hd__and3_1
X_09199_ _13540_/Q _09206_/B VGND VGND VPWR VPWR _09210_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11230_ _10944_/A _11227_/Y _11229_/Y _10929_/A VGND VGND VPWR VPWR _11231_/B sky130_fd_sc_hd__a211o_1
XFILLER_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11161_ _11161_/A VGND VGND VPWR VPWR _11161_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10112_ _10121_/S VGND VGND VPWR VPWR _10119_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_96_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11092_ _11092_/A VGND VGND VPWR VPWR _11092_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10043_ _10043_/A VGND VGND VPWR VPWR _13947_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_152_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold62 hold62/A VGND VGND VPWR VPWR hold62/X sky130_fd_sc_hd__clkbuf_2
Xhold73 hold73/A VGND VGND VPWR VPWR hold73/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_152_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold84 hold84/A VGND VGND VPWR VPWR hold84/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold95 hold95/A VGND VGND VPWR VPWR hold95/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_152_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13802_ _13945_/CLK _13802_/D VGND VGND VPWR VPWR _13802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11994_ _14518_/Q VGND VGND VPWR VPWR _11994_/X sky130_fd_sc_hd__buf_2
XFILLER_44_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13733_ _13805_/CLK hold291/X VGND VGND VPWR VPWR _13733_/Q sky130_fd_sc_hd__dfxtp_1
X_10945_ _11166_/A VGND VGND VPWR VPWR _11224_/A sky130_fd_sc_hd__buf_2
XFILLER_32_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13664_ _13666_/CLK _13664_/D VGND VGND VPWR VPWR _13664_/Q sky130_fd_sc_hd__dfxtp_1
X_10876_ _10876_/A VGND VGND VPWR VPWR _10885_/B sky130_fd_sc_hd__clkbuf_1
X_12615_ _12604_/C _12614_/Y _12580_/X VGND VGND VPWR VPWR _14735_/D sky130_fd_sc_hd__o21a_1
XFILLER_31_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13595_ _13596_/CLK _13595_/D repeater56/X VGND VGND VPWR VPWR _13595_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12546_ _11329_/X _14718_/Q _12554_/S VGND VGND VPWR VPWR _12547_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12477_ _12477_/A VGND VGND VPWR VPWR _14669_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_4 _12261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14216_ _14440_/CLK _14216_/D VGND VGND VPWR VPWR _14216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11428_ _11428_/A VGND VGND VPWR VPWR _13805_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14147_ _14294_/CLK hold184/X VGND VGND VPWR VPWR hold400/A sky130_fd_sc_hd__dfxtp_1
X_11359_ _12016_/A VGND VGND VPWR VPWR _11359_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14078_ _14610_/CLK hold299/X VGND VGND VPWR VPWR hold317/A sky130_fd_sc_hd__dfxtp_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05920_ _13734_/Q _13735_/Q _13736_/Q _05920_/D VGND VGND VPWR VPWR _05921_/D sky130_fd_sc_hd__or4_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ _14108_/CLK _13029_/D repeater59/X VGND VGND VPWR VPWR _13029_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_66_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08570_ _08570_/A VGND VGND VPWR VPWR _08577_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_54_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07521_ _13153_/Q _09228_/B VGND VGND VPWR VPWR _07522_/B sky130_fd_sc_hd__nor2_1
XFILLER_35_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07452_ _07452_/A _07452_/B VGND VGND VPWR VPWR _07454_/C sky130_fd_sc_hd__or2_2
XFILLER_34_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06403_ _06429_/A VGND VGND VPWR VPWR _06471_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_07383_ _07416_/B _07383_/B VGND VGND VPWR VPWR _07383_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_22_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09122_ _09134_/C _09122_/B VGND VGND VPWR VPWR _09122_/X sky130_fd_sc_hd__or2_1
XFILLER_148_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06334_ _06334_/A VGND VGND VPWR VPWR _14402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09053_ _13700_/D VGND VGND VPWR VPWR _09644_/A sky130_fd_sc_hd__buf_2
X_06265_ _06265_/A VGND VGND VPWR VPWR _13977_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08004_ _08013_/A _08013_/B VGND VGND VPWR VPWR _08004_/Y sky130_fd_sc_hd__nor2_1
Xhold510 hold510/A VGND VGND VPWR VPWR hold510/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_06196_ _14420_/Q _14418_/Q _10194_/A VGND VGND VPWR VPWR _06196_/X sky130_fd_sc_hd__mux2_1
Xhold521 hold521/A VGND VGND VPWR VPWR hold521/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_131_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09955_ _13501_/Q _13690_/Q _09957_/S VGND VGND VPWR VPWR _09956_/A sky130_fd_sc_hd__mux2_1
X_08906_ _08927_/A _08978_/B _08978_/D _08907_/A VGND VGND VPWR VPWR _08908_/A sky130_fd_sc_hd__a22oi_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _09886_/A VGND VGND VPWR VPWR _09893_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08837_ _08847_/A _08837_/B VGND VGND VPWR VPWR _08846_/B sky130_fd_sc_hd__xnor2_1
XFILLER_85_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _08770_/B _08768_/B VGND VGND VPWR VPWR _08768_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_72_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07719_ _07684_/Y _07718_/Y _07781_/S VGND VGND VPWR VPWR _07720_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ _13453_/Q _08730_/B VGND VGND VPWR VPWR _08709_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10730_ _10730_/A VGND VGND VPWR VPWR _12942_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10661_ _10666_/C _10673_/B _10661_/C VGND VGND VPWR VPWR _10662_/A sky130_fd_sc_hd__and3b_1
XFILLER_41_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12400_ input17/X _12402_/B _12400_/C VGND VGND VPWR VPWR _12401_/A sky130_fd_sc_hd__and3_1
X_13380_ _14333_/CLK _13380_/D _12609_/A VGND VGND VPWR VPWR _13380_/Q sky130_fd_sc_hd__dfrtp_1
X_10592_ _14583_/Q _10592_/B VGND VGND VPWR VPWR _13746_/D sky130_fd_sc_hd__xor2_1
X_12331_ _12331_/A VGND VGND VPWR VPWR _14580_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12262_ _11329_/X _14546_/Q _12270_/S VGND VGND VPWR VPWR _12263_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11213_ _11207_/X _11210_/X _11212_/X _11157_/X VGND VGND VPWR VPWR _11213_/X sky130_fd_sc_hd__o211a_1
X_14001_ _14725_/CLK _14001_/D VGND VGND VPWR VPWR _14001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12193_ _12193_/A VGND VGND VPWR VPWR _14507_/D sky130_fd_sc_hd__clkbuf_1
Xoutput30 _13318_/Q VGND VGND VPWR VPWR data_o[0] sky130_fd_sc_hd__buf_2
Xoutput41 _13319_/Q VGND VGND VPWR VPWR data_o[1] sky130_fd_sc_hd__buf_2
Xoutput52 _13326_/Q VGND VGND VPWR VPWR data_o[8] sky130_fd_sc_hd__buf_2
X_11144_ _11144_/A VGND VGND VPWR VPWR _11144_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11075_ _11106_/A _11075_/B VGND VGND VPWR VPWR _11075_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10026_ _10606_/C _10024_/X _10032_/S VGND VGND VPWR VPWR _10027_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11977_ _11977_/A VGND VGND VPWR VPWR _14302_/D sky130_fd_sc_hd__clkbuf_1
X_13716_ _13799_/CLK hold335/X VGND VGND VPWR VPWR _13716_/Q sky130_fd_sc_hd__dfxtp_1
X_10928_ _11166_/A VGND VGND VPWR VPWR _10929_/A sky130_fd_sc_hd__clkbuf_2
X_14696_ _14696_/CLK hold311/X VGND VGND VPWR VPWR _14696_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13647_ _14327_/CLK hold357/X VGND VGND VPWR VPWR _13647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10859_ _13147_/Q _10863_/B VGND VGND VPWR VPWR _10860_/A sky130_fd_sc_hd__and2_1
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13578_ _14319_/CLK hold54/X VGND VGND VPWR VPWR _13578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12529_ _12529_/A VGND VGND VPWR VPWR _14710_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06050_ _06046_/X _06047_/X _06057_/A VGND VGND VPWR VPWR _06051_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06952_ _13018_/Q _13019_/Q _13020_/Q _13021_/Q _07988_/B VGND VGND VPWR VPWR _06952_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_113_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09740_ _09726_/A _09726_/B _09723_/A VGND VGND VPWR VPWR _09741_/B sky130_fd_sc_hd__o21a_1
XFILLER_140_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
.ends

