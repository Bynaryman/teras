module teras (VGND,
    VPWR,
    clk,
    rst_n,
    rtr_i,
    rtr_o,
    rts_i,
    rts_o,
    data_i,
    data_o);
 input VGND;
 input VPWR;
 input clk;
 input rst_n;
 input rtr_i;
 output rtr_o;
 input rts_i;
 output rts_o;
 input [31:0] data_i;
 output [31:0] data_o;

 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire clknet_0_clk;
 wire clknet_1_0_0_clk;
 wire clknet_1_1_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_9_clk;
 wire \fifo_inst.WR_DATA[0] ;
 wire \fifo_inst.WR_DATA[10] ;
 wire \fifo_inst.WR_DATA[11] ;
 wire \fifo_inst.WR_DATA[12] ;
 wire \fifo_inst.WR_DATA[13] ;
 wire \fifo_inst.WR_DATA[14] ;
 wire \fifo_inst.WR_DATA[15] ;
 wire \fifo_inst.WR_DATA[1] ;
 wire \fifo_inst.WR_DATA[2] ;
 wire \fifo_inst.WR_DATA[3] ;
 wire \fifo_inst.WR_DATA[4] ;
 wire \fifo_inst.WR_DATA[5] ;
 wire \fifo_inst.WR_DATA[6] ;
 wire \fifo_inst.WR_DATA[7] ;
 wire \fifo_inst.WR_DATA[8] ;
 wire \fifo_inst.WR_DATA[9] ;
 wire \fifo_inst.mem.RD1_ADDR[0] ;
 wire \fifo_inst.mem.RD1_ADDR[1] ;
 wire \fifo_inst.mem.RD1_ADDR[2] ;
 wire \fifo_inst.mem.RD1_ADDR[3] ;
 wire \fifo_inst.mem.WR1_ADDR[0] ;
 wire \fifo_inst.mem.WR1_ADDR[1] ;
 wire \fifo_inst.mem.WR1_ADDR[2] ;
 wire \fifo_inst.mem.WR1_ADDR[3] ;
 wire \fifo_inst.mem.rMemory[0][0] ;
 wire \fifo_inst.mem.rMemory[0][10] ;
 wire \fifo_inst.mem.rMemory[0][11] ;
 wire \fifo_inst.mem.rMemory[0][12] ;
 wire \fifo_inst.mem.rMemory[0][13] ;
 wire \fifo_inst.mem.rMemory[0][14] ;
 wire \fifo_inst.mem.rMemory[0][15] ;
 wire \fifo_inst.mem.rMemory[0][16] ;
 wire \fifo_inst.mem.rMemory[0][17] ;
 wire \fifo_inst.mem.rMemory[0][18] ;
 wire \fifo_inst.mem.rMemory[0][19] ;
 wire \fifo_inst.mem.rMemory[0][1] ;
 wire \fifo_inst.mem.rMemory[0][20] ;
 wire \fifo_inst.mem.rMemory[0][21] ;
 wire \fifo_inst.mem.rMemory[0][22] ;
 wire \fifo_inst.mem.rMemory[0][23] ;
 wire \fifo_inst.mem.rMemory[0][2] ;
 wire \fifo_inst.mem.rMemory[0][3] ;
 wire \fifo_inst.mem.rMemory[0][4] ;
 wire \fifo_inst.mem.rMemory[0][5] ;
 wire \fifo_inst.mem.rMemory[0][6] ;
 wire \fifo_inst.mem.rMemory[0][7] ;
 wire \fifo_inst.mem.rMemory[0][8] ;
 wire \fifo_inst.mem.rMemory[0][9] ;
 wire \fifo_inst.mem.rMemory[10][0] ;
 wire \fifo_inst.mem.rMemory[10][10] ;
 wire \fifo_inst.mem.rMemory[10][11] ;
 wire \fifo_inst.mem.rMemory[10][12] ;
 wire \fifo_inst.mem.rMemory[10][13] ;
 wire \fifo_inst.mem.rMemory[10][14] ;
 wire \fifo_inst.mem.rMemory[10][15] ;
 wire \fifo_inst.mem.rMemory[10][16] ;
 wire \fifo_inst.mem.rMemory[10][17] ;
 wire \fifo_inst.mem.rMemory[10][18] ;
 wire \fifo_inst.mem.rMemory[10][19] ;
 wire \fifo_inst.mem.rMemory[10][1] ;
 wire \fifo_inst.mem.rMemory[10][20] ;
 wire \fifo_inst.mem.rMemory[10][21] ;
 wire \fifo_inst.mem.rMemory[10][22] ;
 wire \fifo_inst.mem.rMemory[10][23] ;
 wire \fifo_inst.mem.rMemory[10][2] ;
 wire \fifo_inst.mem.rMemory[10][3] ;
 wire \fifo_inst.mem.rMemory[10][4] ;
 wire \fifo_inst.mem.rMemory[10][5] ;
 wire \fifo_inst.mem.rMemory[10][6] ;
 wire \fifo_inst.mem.rMemory[10][7] ;
 wire \fifo_inst.mem.rMemory[10][8] ;
 wire \fifo_inst.mem.rMemory[10][9] ;
 wire \fifo_inst.mem.rMemory[11][0] ;
 wire \fifo_inst.mem.rMemory[11][10] ;
 wire \fifo_inst.mem.rMemory[11][11] ;
 wire \fifo_inst.mem.rMemory[11][12] ;
 wire \fifo_inst.mem.rMemory[11][13] ;
 wire \fifo_inst.mem.rMemory[11][14] ;
 wire \fifo_inst.mem.rMemory[11][15] ;
 wire \fifo_inst.mem.rMemory[11][16] ;
 wire \fifo_inst.mem.rMemory[11][17] ;
 wire \fifo_inst.mem.rMemory[11][18] ;
 wire \fifo_inst.mem.rMemory[11][19] ;
 wire \fifo_inst.mem.rMemory[11][1] ;
 wire \fifo_inst.mem.rMemory[11][20] ;
 wire \fifo_inst.mem.rMemory[11][21] ;
 wire \fifo_inst.mem.rMemory[11][22] ;
 wire \fifo_inst.mem.rMemory[11][23] ;
 wire \fifo_inst.mem.rMemory[11][2] ;
 wire \fifo_inst.mem.rMemory[11][3] ;
 wire \fifo_inst.mem.rMemory[11][4] ;
 wire \fifo_inst.mem.rMemory[11][5] ;
 wire \fifo_inst.mem.rMemory[11][6] ;
 wire \fifo_inst.mem.rMemory[11][7] ;
 wire \fifo_inst.mem.rMemory[11][8] ;
 wire \fifo_inst.mem.rMemory[11][9] ;
 wire \fifo_inst.mem.rMemory[12][0] ;
 wire \fifo_inst.mem.rMemory[12][10] ;
 wire \fifo_inst.mem.rMemory[12][11] ;
 wire \fifo_inst.mem.rMemory[12][12] ;
 wire \fifo_inst.mem.rMemory[12][13] ;
 wire \fifo_inst.mem.rMemory[12][14] ;
 wire \fifo_inst.mem.rMemory[12][15] ;
 wire \fifo_inst.mem.rMemory[12][16] ;
 wire \fifo_inst.mem.rMemory[12][17] ;
 wire \fifo_inst.mem.rMemory[12][18] ;
 wire \fifo_inst.mem.rMemory[12][19] ;
 wire \fifo_inst.mem.rMemory[12][1] ;
 wire \fifo_inst.mem.rMemory[12][20] ;
 wire \fifo_inst.mem.rMemory[12][21] ;
 wire \fifo_inst.mem.rMemory[12][22] ;
 wire \fifo_inst.mem.rMemory[12][23] ;
 wire \fifo_inst.mem.rMemory[12][2] ;
 wire \fifo_inst.mem.rMemory[12][3] ;
 wire \fifo_inst.mem.rMemory[12][4] ;
 wire \fifo_inst.mem.rMemory[12][5] ;
 wire \fifo_inst.mem.rMemory[12][6] ;
 wire \fifo_inst.mem.rMemory[12][7] ;
 wire \fifo_inst.mem.rMemory[12][8] ;
 wire \fifo_inst.mem.rMemory[12][9] ;
 wire \fifo_inst.mem.rMemory[13][0] ;
 wire \fifo_inst.mem.rMemory[13][10] ;
 wire \fifo_inst.mem.rMemory[13][11] ;
 wire \fifo_inst.mem.rMemory[13][12] ;
 wire \fifo_inst.mem.rMemory[13][13] ;
 wire \fifo_inst.mem.rMemory[13][14] ;
 wire \fifo_inst.mem.rMemory[13][15] ;
 wire \fifo_inst.mem.rMemory[13][16] ;
 wire \fifo_inst.mem.rMemory[13][17] ;
 wire \fifo_inst.mem.rMemory[13][18] ;
 wire \fifo_inst.mem.rMemory[13][19] ;
 wire \fifo_inst.mem.rMemory[13][1] ;
 wire \fifo_inst.mem.rMemory[13][20] ;
 wire \fifo_inst.mem.rMemory[13][21] ;
 wire \fifo_inst.mem.rMemory[13][22] ;
 wire \fifo_inst.mem.rMemory[13][23] ;
 wire \fifo_inst.mem.rMemory[13][2] ;
 wire \fifo_inst.mem.rMemory[13][3] ;
 wire \fifo_inst.mem.rMemory[13][4] ;
 wire \fifo_inst.mem.rMemory[13][5] ;
 wire \fifo_inst.mem.rMemory[13][6] ;
 wire \fifo_inst.mem.rMemory[13][7] ;
 wire \fifo_inst.mem.rMemory[13][8] ;
 wire \fifo_inst.mem.rMemory[13][9] ;
 wire \fifo_inst.mem.rMemory[14][0] ;
 wire \fifo_inst.mem.rMemory[14][10] ;
 wire \fifo_inst.mem.rMemory[14][11] ;
 wire \fifo_inst.mem.rMemory[14][12] ;
 wire \fifo_inst.mem.rMemory[14][13] ;
 wire \fifo_inst.mem.rMemory[14][14] ;
 wire \fifo_inst.mem.rMemory[14][15] ;
 wire \fifo_inst.mem.rMemory[14][16] ;
 wire \fifo_inst.mem.rMemory[14][17] ;
 wire \fifo_inst.mem.rMemory[14][18] ;
 wire \fifo_inst.mem.rMemory[14][19] ;
 wire \fifo_inst.mem.rMemory[14][1] ;
 wire \fifo_inst.mem.rMemory[14][20] ;
 wire \fifo_inst.mem.rMemory[14][21] ;
 wire \fifo_inst.mem.rMemory[14][22] ;
 wire \fifo_inst.mem.rMemory[14][23] ;
 wire \fifo_inst.mem.rMemory[14][2] ;
 wire \fifo_inst.mem.rMemory[14][3] ;
 wire \fifo_inst.mem.rMemory[14][4] ;
 wire \fifo_inst.mem.rMemory[14][5] ;
 wire \fifo_inst.mem.rMemory[14][6] ;
 wire \fifo_inst.mem.rMemory[14][7] ;
 wire \fifo_inst.mem.rMemory[14][8] ;
 wire \fifo_inst.mem.rMemory[14][9] ;
 wire \fifo_inst.mem.rMemory[15][0] ;
 wire \fifo_inst.mem.rMemory[15][10] ;
 wire \fifo_inst.mem.rMemory[15][11] ;
 wire \fifo_inst.mem.rMemory[15][12] ;
 wire \fifo_inst.mem.rMemory[15][13] ;
 wire \fifo_inst.mem.rMemory[15][14] ;
 wire \fifo_inst.mem.rMemory[15][15] ;
 wire \fifo_inst.mem.rMemory[15][16] ;
 wire \fifo_inst.mem.rMemory[15][17] ;
 wire \fifo_inst.mem.rMemory[15][18] ;
 wire \fifo_inst.mem.rMemory[15][19] ;
 wire \fifo_inst.mem.rMemory[15][1] ;
 wire \fifo_inst.mem.rMemory[15][20] ;
 wire \fifo_inst.mem.rMemory[15][21] ;
 wire \fifo_inst.mem.rMemory[15][22] ;
 wire \fifo_inst.mem.rMemory[15][23] ;
 wire \fifo_inst.mem.rMemory[15][2] ;
 wire \fifo_inst.mem.rMemory[15][3] ;
 wire \fifo_inst.mem.rMemory[15][4] ;
 wire \fifo_inst.mem.rMemory[15][5] ;
 wire \fifo_inst.mem.rMemory[15][6] ;
 wire \fifo_inst.mem.rMemory[15][7] ;
 wire \fifo_inst.mem.rMemory[15][8] ;
 wire \fifo_inst.mem.rMemory[15][9] ;
 wire \fifo_inst.mem.rMemory[1][0] ;
 wire \fifo_inst.mem.rMemory[1][10] ;
 wire \fifo_inst.mem.rMemory[1][11] ;
 wire \fifo_inst.mem.rMemory[1][12] ;
 wire \fifo_inst.mem.rMemory[1][13] ;
 wire \fifo_inst.mem.rMemory[1][14] ;
 wire \fifo_inst.mem.rMemory[1][15] ;
 wire \fifo_inst.mem.rMemory[1][16] ;
 wire \fifo_inst.mem.rMemory[1][17] ;
 wire \fifo_inst.mem.rMemory[1][18] ;
 wire \fifo_inst.mem.rMemory[1][19] ;
 wire \fifo_inst.mem.rMemory[1][1] ;
 wire \fifo_inst.mem.rMemory[1][20] ;
 wire \fifo_inst.mem.rMemory[1][21] ;
 wire \fifo_inst.mem.rMemory[1][22] ;
 wire \fifo_inst.mem.rMemory[1][23] ;
 wire \fifo_inst.mem.rMemory[1][2] ;
 wire \fifo_inst.mem.rMemory[1][3] ;
 wire \fifo_inst.mem.rMemory[1][4] ;
 wire \fifo_inst.mem.rMemory[1][5] ;
 wire \fifo_inst.mem.rMemory[1][6] ;
 wire \fifo_inst.mem.rMemory[1][7] ;
 wire \fifo_inst.mem.rMemory[1][8] ;
 wire \fifo_inst.mem.rMemory[1][9] ;
 wire \fifo_inst.mem.rMemory[2][0] ;
 wire \fifo_inst.mem.rMemory[2][10] ;
 wire \fifo_inst.mem.rMemory[2][11] ;
 wire \fifo_inst.mem.rMemory[2][12] ;
 wire \fifo_inst.mem.rMemory[2][13] ;
 wire \fifo_inst.mem.rMemory[2][14] ;
 wire \fifo_inst.mem.rMemory[2][15] ;
 wire \fifo_inst.mem.rMemory[2][16] ;
 wire \fifo_inst.mem.rMemory[2][17] ;
 wire \fifo_inst.mem.rMemory[2][18] ;
 wire \fifo_inst.mem.rMemory[2][19] ;
 wire \fifo_inst.mem.rMemory[2][1] ;
 wire \fifo_inst.mem.rMemory[2][20] ;
 wire \fifo_inst.mem.rMemory[2][21] ;
 wire \fifo_inst.mem.rMemory[2][22] ;
 wire \fifo_inst.mem.rMemory[2][23] ;
 wire \fifo_inst.mem.rMemory[2][2] ;
 wire \fifo_inst.mem.rMemory[2][3] ;
 wire \fifo_inst.mem.rMemory[2][4] ;
 wire \fifo_inst.mem.rMemory[2][5] ;
 wire \fifo_inst.mem.rMemory[2][6] ;
 wire \fifo_inst.mem.rMemory[2][7] ;
 wire \fifo_inst.mem.rMemory[2][8] ;
 wire \fifo_inst.mem.rMemory[2][9] ;
 wire \fifo_inst.mem.rMemory[3][0] ;
 wire \fifo_inst.mem.rMemory[3][10] ;
 wire \fifo_inst.mem.rMemory[3][11] ;
 wire \fifo_inst.mem.rMemory[3][12] ;
 wire \fifo_inst.mem.rMemory[3][13] ;
 wire \fifo_inst.mem.rMemory[3][14] ;
 wire \fifo_inst.mem.rMemory[3][15] ;
 wire \fifo_inst.mem.rMemory[3][16] ;
 wire \fifo_inst.mem.rMemory[3][17] ;
 wire \fifo_inst.mem.rMemory[3][18] ;
 wire \fifo_inst.mem.rMemory[3][19] ;
 wire \fifo_inst.mem.rMemory[3][1] ;
 wire \fifo_inst.mem.rMemory[3][20] ;
 wire \fifo_inst.mem.rMemory[3][21] ;
 wire \fifo_inst.mem.rMemory[3][22] ;
 wire \fifo_inst.mem.rMemory[3][23] ;
 wire \fifo_inst.mem.rMemory[3][2] ;
 wire \fifo_inst.mem.rMemory[3][3] ;
 wire \fifo_inst.mem.rMemory[3][4] ;
 wire \fifo_inst.mem.rMemory[3][5] ;
 wire \fifo_inst.mem.rMemory[3][6] ;
 wire \fifo_inst.mem.rMemory[3][7] ;
 wire \fifo_inst.mem.rMemory[3][8] ;
 wire \fifo_inst.mem.rMemory[3][9] ;
 wire \fifo_inst.mem.rMemory[4][0] ;
 wire \fifo_inst.mem.rMemory[4][10] ;
 wire \fifo_inst.mem.rMemory[4][11] ;
 wire \fifo_inst.mem.rMemory[4][12] ;
 wire \fifo_inst.mem.rMemory[4][13] ;
 wire \fifo_inst.mem.rMemory[4][14] ;
 wire \fifo_inst.mem.rMemory[4][15] ;
 wire \fifo_inst.mem.rMemory[4][16] ;
 wire \fifo_inst.mem.rMemory[4][17] ;
 wire \fifo_inst.mem.rMemory[4][18] ;
 wire \fifo_inst.mem.rMemory[4][19] ;
 wire \fifo_inst.mem.rMemory[4][1] ;
 wire \fifo_inst.mem.rMemory[4][20] ;
 wire \fifo_inst.mem.rMemory[4][21] ;
 wire \fifo_inst.mem.rMemory[4][22] ;
 wire \fifo_inst.mem.rMemory[4][23] ;
 wire \fifo_inst.mem.rMemory[4][2] ;
 wire \fifo_inst.mem.rMemory[4][3] ;
 wire \fifo_inst.mem.rMemory[4][4] ;
 wire \fifo_inst.mem.rMemory[4][5] ;
 wire \fifo_inst.mem.rMemory[4][6] ;
 wire \fifo_inst.mem.rMemory[4][7] ;
 wire \fifo_inst.mem.rMemory[4][8] ;
 wire \fifo_inst.mem.rMemory[4][9] ;
 wire \fifo_inst.mem.rMemory[5][0] ;
 wire \fifo_inst.mem.rMemory[5][10] ;
 wire \fifo_inst.mem.rMemory[5][11] ;
 wire \fifo_inst.mem.rMemory[5][12] ;
 wire \fifo_inst.mem.rMemory[5][13] ;
 wire \fifo_inst.mem.rMemory[5][14] ;
 wire \fifo_inst.mem.rMemory[5][15] ;
 wire \fifo_inst.mem.rMemory[5][16] ;
 wire \fifo_inst.mem.rMemory[5][17] ;
 wire \fifo_inst.mem.rMemory[5][18] ;
 wire \fifo_inst.mem.rMemory[5][19] ;
 wire \fifo_inst.mem.rMemory[5][1] ;
 wire \fifo_inst.mem.rMemory[5][20] ;
 wire \fifo_inst.mem.rMemory[5][21] ;
 wire \fifo_inst.mem.rMemory[5][22] ;
 wire \fifo_inst.mem.rMemory[5][23] ;
 wire \fifo_inst.mem.rMemory[5][2] ;
 wire \fifo_inst.mem.rMemory[5][3] ;
 wire \fifo_inst.mem.rMemory[5][4] ;
 wire \fifo_inst.mem.rMemory[5][5] ;
 wire \fifo_inst.mem.rMemory[5][6] ;
 wire \fifo_inst.mem.rMemory[5][7] ;
 wire \fifo_inst.mem.rMemory[5][8] ;
 wire \fifo_inst.mem.rMemory[5][9] ;
 wire \fifo_inst.mem.rMemory[6][0] ;
 wire \fifo_inst.mem.rMemory[6][10] ;
 wire \fifo_inst.mem.rMemory[6][11] ;
 wire \fifo_inst.mem.rMemory[6][12] ;
 wire \fifo_inst.mem.rMemory[6][13] ;
 wire \fifo_inst.mem.rMemory[6][14] ;
 wire \fifo_inst.mem.rMemory[6][15] ;
 wire \fifo_inst.mem.rMemory[6][16] ;
 wire \fifo_inst.mem.rMemory[6][17] ;
 wire \fifo_inst.mem.rMemory[6][18] ;
 wire \fifo_inst.mem.rMemory[6][19] ;
 wire \fifo_inst.mem.rMemory[6][1] ;
 wire \fifo_inst.mem.rMemory[6][20] ;
 wire \fifo_inst.mem.rMemory[6][21] ;
 wire \fifo_inst.mem.rMemory[6][22] ;
 wire \fifo_inst.mem.rMemory[6][23] ;
 wire \fifo_inst.mem.rMemory[6][2] ;
 wire \fifo_inst.mem.rMemory[6][3] ;
 wire \fifo_inst.mem.rMemory[6][4] ;
 wire \fifo_inst.mem.rMemory[6][5] ;
 wire \fifo_inst.mem.rMemory[6][6] ;
 wire \fifo_inst.mem.rMemory[6][7] ;
 wire \fifo_inst.mem.rMemory[6][8] ;
 wire \fifo_inst.mem.rMemory[6][9] ;
 wire \fifo_inst.mem.rMemory[7][0] ;
 wire \fifo_inst.mem.rMemory[7][10] ;
 wire \fifo_inst.mem.rMemory[7][11] ;
 wire \fifo_inst.mem.rMemory[7][12] ;
 wire \fifo_inst.mem.rMemory[7][13] ;
 wire \fifo_inst.mem.rMemory[7][14] ;
 wire \fifo_inst.mem.rMemory[7][15] ;
 wire \fifo_inst.mem.rMemory[7][16] ;
 wire \fifo_inst.mem.rMemory[7][17] ;
 wire \fifo_inst.mem.rMemory[7][18] ;
 wire \fifo_inst.mem.rMemory[7][19] ;
 wire \fifo_inst.mem.rMemory[7][1] ;
 wire \fifo_inst.mem.rMemory[7][20] ;
 wire \fifo_inst.mem.rMemory[7][21] ;
 wire \fifo_inst.mem.rMemory[7][22] ;
 wire \fifo_inst.mem.rMemory[7][23] ;
 wire \fifo_inst.mem.rMemory[7][2] ;
 wire \fifo_inst.mem.rMemory[7][3] ;
 wire \fifo_inst.mem.rMemory[7][4] ;
 wire \fifo_inst.mem.rMemory[7][5] ;
 wire \fifo_inst.mem.rMemory[7][6] ;
 wire \fifo_inst.mem.rMemory[7][7] ;
 wire \fifo_inst.mem.rMemory[7][8] ;
 wire \fifo_inst.mem.rMemory[7][9] ;
 wire \fifo_inst.mem.rMemory[8][0] ;
 wire \fifo_inst.mem.rMemory[8][10] ;
 wire \fifo_inst.mem.rMemory[8][11] ;
 wire \fifo_inst.mem.rMemory[8][12] ;
 wire \fifo_inst.mem.rMemory[8][13] ;
 wire \fifo_inst.mem.rMemory[8][14] ;
 wire \fifo_inst.mem.rMemory[8][15] ;
 wire \fifo_inst.mem.rMemory[8][16] ;
 wire \fifo_inst.mem.rMemory[8][17] ;
 wire \fifo_inst.mem.rMemory[8][18] ;
 wire \fifo_inst.mem.rMemory[8][19] ;
 wire \fifo_inst.mem.rMemory[8][1] ;
 wire \fifo_inst.mem.rMemory[8][20] ;
 wire \fifo_inst.mem.rMemory[8][21] ;
 wire \fifo_inst.mem.rMemory[8][22] ;
 wire \fifo_inst.mem.rMemory[8][23] ;
 wire \fifo_inst.mem.rMemory[8][2] ;
 wire \fifo_inst.mem.rMemory[8][3] ;
 wire \fifo_inst.mem.rMemory[8][4] ;
 wire \fifo_inst.mem.rMemory[8][5] ;
 wire \fifo_inst.mem.rMemory[8][6] ;
 wire \fifo_inst.mem.rMemory[8][7] ;
 wire \fifo_inst.mem.rMemory[8][8] ;
 wire \fifo_inst.mem.rMemory[8][9] ;
 wire \fifo_inst.mem.rMemory[9][0] ;
 wire \fifo_inst.mem.rMemory[9][10] ;
 wire \fifo_inst.mem.rMemory[9][11] ;
 wire \fifo_inst.mem.rMemory[9][12] ;
 wire \fifo_inst.mem.rMemory[9][13] ;
 wire \fifo_inst.mem.rMemory[9][14] ;
 wire \fifo_inst.mem.rMemory[9][15] ;
 wire \fifo_inst.mem.rMemory[9][16] ;
 wire \fifo_inst.mem.rMemory[9][17] ;
 wire \fifo_inst.mem.rMemory[9][18] ;
 wire \fifo_inst.mem.rMemory[9][19] ;
 wire \fifo_inst.mem.rMemory[9][1] ;
 wire \fifo_inst.mem.rMemory[9][20] ;
 wire \fifo_inst.mem.rMemory[9][21] ;
 wire \fifo_inst.mem.rMemory[9][22] ;
 wire \fifo_inst.mem.rMemory[9][23] ;
 wire \fifo_inst.mem.rMemory[9][2] ;
 wire \fifo_inst.mem.rMemory[9][3] ;
 wire \fifo_inst.mem.rMemory[9][4] ;
 wire \fifo_inst.mem.rMemory[9][5] ;
 wire \fifo_inst.mem.rMemory[9][6] ;
 wire \fifo_inst.mem.rMemory[9][7] ;
 wire \fifo_inst.mem.rMemory[9][8] ;
 wire \fifo_inst.mem.rMemory[9][9] ;
 wire \fifo_inst.rEmpty ;
 wire \fifo_inst.rFull ;
 wire \fifo_inst.rRdPtrPlus1[0] ;
 wire \fifo_inst.rRdPtrPlus1[1] ;
 wire \fifo_inst.rRdPtrPlus1[2] ;
 wire \fifo_inst.rRdPtrPlus1[3] ;
 wire \fifo_inst.rRdPtrPlus1[4] ;
 wire \fifo_inst.rRdPtr[4] ;
 wire \fifo_inst.rWrPtrPlus1[0] ;
 wire \fifo_inst.rWrPtrPlus1[1] ;
 wire \fifo_inst.rWrPtrPlus1[2] ;
 wire \fifo_inst.rWrPtrPlus1[3] ;
 wire \fifo_inst.rWrPtrPlus1[4] ;
 wire \fifo_inst.rWrPtr[4] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net8;
 wire net9;
 wire \sa_inst.EOB_Q_o ;
 wire \sa_inst._00_[0] ;
 wire \sa_inst._00_[1] ;
 wire \sa_inst._00_[2] ;
 wire \sa_inst._00_[3] ;
 wire \sa_inst._00_[4] ;
 wire \sa_inst._00_[5] ;
 wire \sa_inst._00_[6] ;
 wire \sa_inst._00_[7] ;
 wire \sa_inst._01_ ;
 wire \sa_inst._02_[0] ;
 wire \sa_inst._02_[1] ;
 wire \sa_inst._02_[2] ;
 wire \sa_inst._02_[3] ;
 wire \sa_inst._02_[4] ;
 wire \sa_inst._02_[5] ;
 wire \sa_inst._02_[6] ;
 wire \sa_inst._02_[7] ;
 wire \sa_inst._05_[0] ;
 wire \sa_inst._05_[10] ;
 wire \sa_inst._05_[11] ;
 wire \sa_inst._05_[1] ;
 wire \sa_inst._05_[2] ;
 wire \sa_inst._05_[3] ;
 wire \sa_inst._05_[4] ;
 wire \sa_inst._05_[5] ;
 wire \sa_inst._05_[6] ;
 wire \sa_inst._05_[7] ;
 wire \sa_inst._05_[8] ;
 wire \sa_inst._05_[9] ;
 wire \sa_inst._06_[0] ;
 wire \sa_inst._06_[10] ;
 wire \sa_inst._06_[11] ;
 wire \sa_inst._06_[1] ;
 wire \sa_inst._06_[2] ;
 wire \sa_inst._06_[3] ;
 wire \sa_inst._06_[4] ;
 wire \sa_inst._06_[5] ;
 wire \sa_inst._06_[6] ;
 wire \sa_inst._06_[7] ;
 wire \sa_inst._06_[8] ;
 wire \sa_inst._06_[9] ;
 wire \sa_inst._07_[0] ;
 wire \sa_inst._07_[10] ;
 wire \sa_inst._07_[11] ;
 wire \sa_inst._07_[1] ;
 wire \sa_inst._07_[2] ;
 wire \sa_inst._07_[3] ;
 wire \sa_inst._07_[4] ;
 wire \sa_inst._07_[5] ;
 wire \sa_inst._07_[6] ;
 wire \sa_inst._07_[7] ;
 wire \sa_inst._07_[8] ;
 wire \sa_inst._07_[9] ;
 wire \sa_inst._11_[0] ;
 wire \sa_inst._11_[1] ;
 wire \sa_inst._11_[2] ;
 wire \sa_inst._11_[3] ;
 wire \sa_inst._11_[4] ;
 wire \sa_inst._11_[5] ;
 wire \sa_inst._11_[6] ;
 wire \sa_inst._11_[7] ;
 wire \sa_inst._12_[0] ;
 wire \sa_inst._12_[10] ;
 wire \sa_inst._12_[11] ;
 wire \sa_inst._12_[12] ;
 wire \sa_inst._12_[13] ;
 wire \sa_inst._12_[14] ;
 wire \sa_inst._12_[15] ;
 wire \sa_inst._12_[16] ;
 wire \sa_inst._12_[17] ;
 wire \sa_inst._12_[18] ;
 wire \sa_inst._12_[19] ;
 wire \sa_inst._12_[1] ;
 wire \sa_inst._12_[20] ;
 wire \sa_inst._12_[21] ;
 wire \sa_inst._12_[22] ;
 wire \sa_inst._12_[23] ;
 wire \sa_inst._12_[24] ;
 wire \sa_inst._12_[25] ;
 wire \sa_inst._12_[26] ;
 wire \sa_inst._12_[27] ;
 wire \sa_inst._12_[28] ;
 wire \sa_inst._12_[29] ;
 wire \sa_inst._12_[2] ;
 wire \sa_inst._12_[30] ;
 wire \sa_inst._12_[31] ;
 wire \sa_inst._12_[32] ;
 wire \sa_inst._12_[33] ;
 wire \sa_inst._12_[34] ;
 wire \sa_inst._12_[35] ;
 wire \sa_inst._12_[36] ;
 wire \sa_inst._12_[37] ;
 wire \sa_inst._12_[38] ;
 wire \sa_inst._12_[39] ;
 wire \sa_inst._12_[3] ;
 wire \sa_inst._12_[40] ;
 wire \sa_inst._12_[41] ;
 wire \sa_inst._12_[42] ;
 wire \sa_inst._12_[43] ;
 wire \sa_inst._12_[44] ;
 wire \sa_inst._12_[45] ;
 wire \sa_inst._12_[46] ;
 wire \sa_inst._12_[47] ;
 wire \sa_inst._12_[48] ;
 wire \sa_inst._12_[49] ;
 wire \sa_inst._12_[4] ;
 wire \sa_inst._12_[50] ;
 wire \sa_inst._12_[51] ;
 wire \sa_inst._12_[52] ;
 wire \sa_inst._12_[53] ;
 wire \sa_inst._12_[54] ;
 wire \sa_inst._12_[55] ;
 wire \sa_inst._12_[56] ;
 wire \sa_inst._12_[57] ;
 wire \sa_inst._12_[58] ;
 wire \sa_inst._12_[59] ;
 wire \sa_inst._12_[5] ;
 wire \sa_inst._12_[60] ;
 wire \sa_inst._12_[61] ;
 wire \sa_inst._12_[62] ;
 wire \sa_inst._12_[63] ;
 wire \sa_inst._12_[64] ;
 wire \sa_inst._12_[65] ;
 wire \sa_inst._12_[66] ;
 wire \sa_inst._12_[67] ;
 wire \sa_inst._12_[68] ;
 wire \sa_inst._12_[69] ;
 wire \sa_inst._12_[6] ;
 wire \sa_inst._12_[70] ;
 wire \sa_inst._12_[71] ;
 wire \sa_inst._12_[72] ;
 wire \sa_inst._12_[73] ;
 wire \sa_inst._12_[74] ;
 wire \sa_inst._12_[75] ;
 wire \sa_inst._12_[76] ;
 wire \sa_inst._12_[77] ;
 wire \sa_inst._12_[78] ;
 wire \sa_inst._12_[79] ;
 wire \sa_inst._12_[7] ;
 wire \sa_inst._12_[80] ;
 wire \sa_inst._12_[81] ;
 wire \sa_inst._12_[82] ;
 wire \sa_inst._12_[83] ;
 wire \sa_inst._12_[84] ;
 wire \sa_inst._12_[85] ;
 wire \sa_inst._12_[86] ;
 wire \sa_inst._12_[87] ;
 wire \sa_inst._12_[88] ;
 wire \sa_inst._12_[89] ;
 wire \sa_inst._12_[8] ;
 wire \sa_inst._12_[90] ;
 wire \sa_inst._12_[91] ;
 wire \sa_inst._12_[92] ;
 wire \sa_inst._12_[93] ;
 wire \sa_inst._12_[94] ;
 wire \sa_inst._12_[95] ;
 wire \sa_inst._12_[96] ;
 wire \sa_inst._12_[97] ;
 wire \sa_inst._12_[98] ;
 wire \sa_inst._12_[9] ;
 wire \sa_inst._17_[0] ;
 wire \sa_inst._17_[1] ;
 wire \sa_inst._17_[2] ;
 wire \sa_inst._17_[3] ;
 wire \sa_inst._17_[4] ;
 wire \sa_inst._17_[5] ;
 wire \sa_inst._17_[6] ;
 wire \sa_inst._17_[7] ;
 wire \sa_inst._21_ ;
 wire \sa_inst._22_ ;
 wire \sa_inst._23_ ;
 wire \sa_inst.arith_in_col_0[6] ;
 wire \sa_inst.arith_in_col_0[7] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._00_ ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._05_ ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._07_ ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._12_[1] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._12_[2] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._12_[3] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._12_[4] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._14_[0] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._15_[0] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._15_[1] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._15_[2] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._15_[3] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._17_ ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._19_ ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._23_[1] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._23_[2] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j._23_[3] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j.lzoc._00_ ;
 wire \sa_inst.cols_a2s3:1.a2s3_j.lzoc._01_ ;
 wire \sa_inst.cols_a2s3:1.a2s3_j.lzoc._08_ ;
 wire \sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[0] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[1] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[2] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[3] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[4] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[5] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j.lzoc._10_ ;
 wire \sa_inst.cols_a2s3:1.a2s3_j.lzoc._11_ ;
 wire \sa_inst.cols_a2s3:1.a2s3_j.lzoc._14_[4] ;
 wire \sa_inst.cols_a2s3:1.a2s3_j.lzoc._14_[5] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j.43$func$/openlane/designs/teras/src/arith_to_s3.v:95$95.$result[0] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j._00_ ;
 wire \sa_inst.cols_a2s3:2.a2s3_j._05_ ;
 wire \sa_inst.cols_a2s3:2.a2s3_j._07_ ;
 wire \sa_inst.cols_a2s3:2.a2s3_j._12_[1] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j._12_[2] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j._12_[3] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j._12_[4] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j._15_[0] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j._15_[1] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j._15_[2] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j._15_[3] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j._17_ ;
 wire \sa_inst.cols_a2s3:2.a2s3_j._19_ ;
 wire \sa_inst.cols_a2s3:2.a2s3_j._23_[1] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j._23_[2] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j._23_[3] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j.lzoc._00_ ;
 wire \sa_inst.cols_a2s3:2.a2s3_j.lzoc._01_ ;
 wire \sa_inst.cols_a2s3:2.a2s3_j.lzoc._08_ ;
 wire \sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[0] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[1] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[2] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[3] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[4] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[5] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j.lzoc._10_ ;
 wire \sa_inst.cols_a2s3:2.a2s3_j.lzoc._11_ ;
 wire \sa_inst.cols_a2s3:2.a2s3_j.lzoc._14_[4] ;
 wire \sa_inst.cols_a2s3:2.a2s3_j.lzoc._14_[5] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j.43$func$/openlane/designs/teras/src/arith_to_s3.v:95$95.$result[0] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j._00_ ;
 wire \sa_inst.cols_a2s3:3.a2s3_j._05_ ;
 wire \sa_inst.cols_a2s3:3.a2s3_j._07_ ;
 wire \sa_inst.cols_a2s3:3.a2s3_j._12_[1] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j._12_[2] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j._12_[3] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j._12_[4] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j._15_[0] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j._15_[1] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j._15_[2] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j._15_[3] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j._17_ ;
 wire \sa_inst.cols_a2s3:3.a2s3_j._19_ ;
 wire \sa_inst.cols_a2s3:3.a2s3_j._23_[1] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j._23_[2] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j._23_[3] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j.lzoc._00_ ;
 wire \sa_inst.cols_a2s3:3.a2s3_j.lzoc._01_ ;
 wire \sa_inst.cols_a2s3:3.a2s3_j.lzoc._08_ ;
 wire \sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[0] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[1] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[2] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[3] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[4] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[5] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j.lzoc._10_ ;
 wire \sa_inst.cols_a2s3:3.a2s3_j.lzoc._11_ ;
 wire \sa_inst.cols_a2s3:3.a2s3_j.lzoc._14_[4] ;
 wire \sa_inst.cols_a2s3:3.a2s3_j.lzoc._14_[5] ;
 wire \sa_inst.cols_l2a:1.l2a_i._00_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._01_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._02_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i._02_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i._02_[2] ;
 wire \sa_inst.cols_l2a:1.l2a_i._02_[3] ;
 wire \sa_inst.cols_l2a:1.l2a_i._02_[4] ;
 wire \sa_inst.cols_l2a:1.l2a_i._02_[5] ;
 wire \sa_inst.cols_l2a:1.l2a_i._03_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i._04_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i._05_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i._05_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i._05_[2] ;
 wire \sa_inst.cols_l2a:1.l2a_i._05_[3] ;
 wire \sa_inst.cols_l2a:1.l2a_i._06_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._07_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i._07_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i._07_[2] ;
 wire \sa_inst.cols_l2a:1.l2a_i._07_[3] ;
 wire \sa_inst.cols_l2a:1.l2a_i._07_[4] ;
 wire \sa_inst.cols_l2a:1.l2a_i._07_[5] ;
 wire \sa_inst.cols_l2a:1.l2a_i._07_[6] ;
 wire \sa_inst.cols_l2a:1.l2a_i._08_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i._08_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i._08_[2] ;
 wire \sa_inst.cols_l2a:1.l2a_i._08_[3] ;
 wire \sa_inst.cols_l2a:1.l2a_i._08_[4] ;
 wire \sa_inst.cols_l2a:1.l2a_i._08_[5] ;
 wire \sa_inst.cols_l2a:1.l2a_i._08_[6] ;
 wire \sa_inst.cols_l2a:1.l2a_i._09_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i._09_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i._09_[2] ;
 wire \sa_inst.cols_l2a:1.l2a_i._09_[3] ;
 wire \sa_inst.cols_l2a:1.l2a_i._09_[4] ;
 wire \sa_inst.cols_l2a:1.l2a_i._09_[5] ;
 wire \sa_inst.cols_l2a:1.l2a_i._09_[6] ;
 wire \sa_inst.cols_l2a:1.l2a_i._11_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._13_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._14_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._15_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._16_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._17_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._18_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._19_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._20_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._21_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._22_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._23_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._24_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._25_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._26_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._27_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._29_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i._29_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i._29_[2] ;
 wire \sa_inst.cols_l2a:1.l2a_i._29_[3] ;
 wire \sa_inst.cols_l2a:1.l2a_i._29_[4] ;
 wire \sa_inst.cols_l2a:1.l2a_i._29_[5] ;
 wire \sa_inst.cols_l2a:1.l2a_i._30_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._31_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i._31_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i._31_[2] ;
 wire \sa_inst.cols_l2a:1.l2a_i._31_[3] ;
 wire \sa_inst.cols_l2a:1.l2a_i._31_[5] ;
 wire \sa_inst.cols_l2a:1.l2a_i._33_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._35_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i._35_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i._35_[2] ;
 wire \sa_inst.cols_l2a:1.l2a_i._35_[3] ;
 wire \sa_inst.cols_l2a:1.l2a_i._37_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._40_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i._40_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i._40_[2] ;
 wire \sa_inst.cols_l2a:1.l2a_i._40_[3] ;
 wire \sa_inst.cols_l2a:1.l2a_i._40_[4] ;
 wire \sa_inst.cols_l2a:1.l2a_i._40_[5] ;
 wire \sa_inst.cols_l2a:1.l2a_i._40_[6] ;
 wire \sa_inst.cols_l2a:1.l2a_i._44_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._46_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._54_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._55_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._56_ ;
 wire \sa_inst.cols_l2a:1.l2a_i._57_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._01_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[10] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[11] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[12] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[13] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[14] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[15] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[16] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[17] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[18] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[19] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[20] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[21] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[22] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[23] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[24] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[25] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[26] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[27] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[28] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[29] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[30] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[8] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[9] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._03_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._05_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._06_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._07_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._08_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._09_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[2] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[3] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[4] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[5] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[6] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[7] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[8] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[9] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._13_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._14_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._15_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._23_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._31_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._33_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[10] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[11] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[12] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[13] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[14] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[15] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[16] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[17] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[18] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[19] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[20] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[21] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[22] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[23] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[24] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[25] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[26] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[27] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[28] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[29] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[30] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[8] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[9] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._42_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._44_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._48_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._50_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._55_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._56_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[2] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[3] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[4] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[5] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[6] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[7] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[8] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[9] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[10] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[11] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[12] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[13] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[14] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[15] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[16] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[17] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[18] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[19] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[20] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[21] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[22] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[23] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[24] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[25] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[26] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[27] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[28] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[29] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[2] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[30] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[31] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[3] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[4] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[5] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[6] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[7] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[8] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[9] ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._67_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._69_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._74_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.lzoc_inst._88_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._00_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._00_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._00_[2] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._04_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._04_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._04_[2] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._04_[3] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._10_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._10_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._11_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._14_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._17_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._18_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._22_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._25_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._25_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._25_[2] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._25_[3] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._26_[0] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._26_[1] ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._27_ ;
 wire \sa_inst.cols_l2a:1.l2a_i.rshift._28_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i._00_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._01_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._02_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i._02_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i._02_[2] ;
 wire \sa_inst.cols_l2a:2.l2a_i._02_[3] ;
 wire \sa_inst.cols_l2a:2.l2a_i._02_[4] ;
 wire \sa_inst.cols_l2a:2.l2a_i._02_[5] ;
 wire \sa_inst.cols_l2a:2.l2a_i._03_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i._04_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i._05_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i._05_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i._05_[2] ;
 wire \sa_inst.cols_l2a:2.l2a_i._05_[3] ;
 wire \sa_inst.cols_l2a:2.l2a_i._06_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._07_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i._07_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i._07_[2] ;
 wire \sa_inst.cols_l2a:2.l2a_i._07_[3] ;
 wire \sa_inst.cols_l2a:2.l2a_i._07_[4] ;
 wire \sa_inst.cols_l2a:2.l2a_i._07_[5] ;
 wire \sa_inst.cols_l2a:2.l2a_i._07_[6] ;
 wire \sa_inst.cols_l2a:2.l2a_i._08_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i._08_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i._08_[2] ;
 wire \sa_inst.cols_l2a:2.l2a_i._08_[3] ;
 wire \sa_inst.cols_l2a:2.l2a_i._08_[4] ;
 wire \sa_inst.cols_l2a:2.l2a_i._08_[5] ;
 wire \sa_inst.cols_l2a:2.l2a_i._08_[6] ;
 wire \sa_inst.cols_l2a:2.l2a_i._09_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i._09_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i._09_[2] ;
 wire \sa_inst.cols_l2a:2.l2a_i._09_[3] ;
 wire \sa_inst.cols_l2a:2.l2a_i._09_[4] ;
 wire \sa_inst.cols_l2a:2.l2a_i._09_[5] ;
 wire \sa_inst.cols_l2a:2.l2a_i._09_[6] ;
 wire \sa_inst.cols_l2a:2.l2a_i._11_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._13_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._14_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._15_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._16_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._17_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._18_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._19_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._20_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._21_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._22_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._23_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._24_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._25_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._26_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._27_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._29_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i._29_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i._29_[2] ;
 wire \sa_inst.cols_l2a:2.l2a_i._29_[3] ;
 wire \sa_inst.cols_l2a:2.l2a_i._29_[4] ;
 wire \sa_inst.cols_l2a:2.l2a_i._29_[5] ;
 wire \sa_inst.cols_l2a:2.l2a_i._30_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._31_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i._31_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i._31_[2] ;
 wire \sa_inst.cols_l2a:2.l2a_i._31_[3] ;
 wire \sa_inst.cols_l2a:2.l2a_i._31_[5] ;
 wire \sa_inst.cols_l2a:2.l2a_i._33_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._35_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i._35_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i._35_[2] ;
 wire \sa_inst.cols_l2a:2.l2a_i._35_[3] ;
 wire \sa_inst.cols_l2a:2.l2a_i._37_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._40_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i._40_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i._40_[2] ;
 wire \sa_inst.cols_l2a:2.l2a_i._40_[3] ;
 wire \sa_inst.cols_l2a:2.l2a_i._40_[4] ;
 wire \sa_inst.cols_l2a:2.l2a_i._40_[5] ;
 wire \sa_inst.cols_l2a:2.l2a_i._40_[6] ;
 wire \sa_inst.cols_l2a:2.l2a_i._44_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._46_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._54_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._55_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._56_ ;
 wire \sa_inst.cols_l2a:2.l2a_i._57_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._01_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[10] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[11] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[12] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[13] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[14] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[15] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[16] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[17] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[18] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[19] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[20] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[21] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[22] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[23] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[24] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[25] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[26] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[27] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[28] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[29] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[30] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[8] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[9] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._03_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._05_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._06_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._07_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._08_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._09_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[2] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[3] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[4] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[5] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[6] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[7] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[8] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[9] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._13_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._14_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._15_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._23_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._31_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._33_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[10] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[11] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[12] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[13] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[14] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[15] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[16] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[17] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[18] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[19] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[20] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[21] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[22] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[23] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[24] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[25] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[26] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[27] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[28] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[29] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[30] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[8] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[9] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._42_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._44_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._48_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._50_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._55_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._56_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[2] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[3] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[4] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[5] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[6] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[7] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[8] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[9] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[10] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[11] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[12] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[13] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[14] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[15] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[16] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[17] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[18] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[19] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[20] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[21] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[22] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[23] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[24] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[25] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[26] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[27] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[28] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[29] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[2] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[30] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[31] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[3] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[4] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[5] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[6] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[7] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[8] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[9] ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._67_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._69_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._74_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.lzoc_inst._88_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._00_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._00_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._00_[2] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._04_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._04_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._04_[2] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._04_[3] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._10_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._10_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._11_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._14_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._17_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._18_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._22_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._25_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._25_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._25_[2] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._25_[3] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._26_[0] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._26_[1] ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._27_ ;
 wire \sa_inst.cols_l2a:2.l2a_i.rshift._28_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i._00_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._01_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._02_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i._02_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i._02_[2] ;
 wire \sa_inst.cols_l2a:3.l2a_i._02_[3] ;
 wire \sa_inst.cols_l2a:3.l2a_i._02_[4] ;
 wire \sa_inst.cols_l2a:3.l2a_i._02_[5] ;
 wire \sa_inst.cols_l2a:3.l2a_i._03_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i._04_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i._05_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i._05_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i._05_[2] ;
 wire \sa_inst.cols_l2a:3.l2a_i._05_[3] ;
 wire \sa_inst.cols_l2a:3.l2a_i._06_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._07_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i._07_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i._07_[2] ;
 wire \sa_inst.cols_l2a:3.l2a_i._07_[3] ;
 wire \sa_inst.cols_l2a:3.l2a_i._07_[4] ;
 wire \sa_inst.cols_l2a:3.l2a_i._07_[5] ;
 wire \sa_inst.cols_l2a:3.l2a_i._07_[6] ;
 wire \sa_inst.cols_l2a:3.l2a_i._08_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i._08_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i._08_[2] ;
 wire \sa_inst.cols_l2a:3.l2a_i._08_[3] ;
 wire \sa_inst.cols_l2a:3.l2a_i._08_[4] ;
 wire \sa_inst.cols_l2a:3.l2a_i._08_[5] ;
 wire \sa_inst.cols_l2a:3.l2a_i._08_[6] ;
 wire \sa_inst.cols_l2a:3.l2a_i._09_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i._09_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i._09_[2] ;
 wire \sa_inst.cols_l2a:3.l2a_i._09_[3] ;
 wire \sa_inst.cols_l2a:3.l2a_i._09_[4] ;
 wire \sa_inst.cols_l2a:3.l2a_i._09_[5] ;
 wire \sa_inst.cols_l2a:3.l2a_i._09_[6] ;
 wire \sa_inst.cols_l2a:3.l2a_i._11_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._13_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._14_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._15_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._16_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._17_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._18_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._19_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._20_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._21_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._22_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._23_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._24_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._25_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._26_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._27_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._29_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i._29_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i._29_[2] ;
 wire \sa_inst.cols_l2a:3.l2a_i._29_[3] ;
 wire \sa_inst.cols_l2a:3.l2a_i._29_[4] ;
 wire \sa_inst.cols_l2a:3.l2a_i._29_[5] ;
 wire \sa_inst.cols_l2a:3.l2a_i._30_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._31_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i._31_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i._31_[2] ;
 wire \sa_inst.cols_l2a:3.l2a_i._31_[3] ;
 wire \sa_inst.cols_l2a:3.l2a_i._31_[5] ;
 wire \sa_inst.cols_l2a:3.l2a_i._33_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._35_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i._35_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i._35_[2] ;
 wire \sa_inst.cols_l2a:3.l2a_i._35_[3] ;
 wire \sa_inst.cols_l2a:3.l2a_i._37_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._40_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i._40_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i._40_[2] ;
 wire \sa_inst.cols_l2a:3.l2a_i._40_[3] ;
 wire \sa_inst.cols_l2a:3.l2a_i._40_[4] ;
 wire \sa_inst.cols_l2a:3.l2a_i._40_[5] ;
 wire \sa_inst.cols_l2a:3.l2a_i._40_[6] ;
 wire \sa_inst.cols_l2a:3.l2a_i._44_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._46_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._54_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._55_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._56_ ;
 wire \sa_inst.cols_l2a:3.l2a_i._57_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._01_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[10] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[11] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[12] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[13] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[14] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[15] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[16] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[17] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[18] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[19] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[20] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[21] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[22] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[23] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[24] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[25] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[26] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[27] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[28] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[29] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[30] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[8] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[9] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._03_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._05_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._06_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._07_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._08_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._09_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[2] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[3] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[4] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[5] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[6] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[7] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[8] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[9] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._13_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._14_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._15_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._23_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._31_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._33_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[10] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[11] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[12] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[13] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[14] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[15] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[16] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[17] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[18] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[19] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[20] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[21] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[22] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[23] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[24] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[25] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[26] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[27] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[28] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[29] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[30] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[8] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[9] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._42_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._44_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._48_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._50_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._55_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._56_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[2] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[3] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[4] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[5] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[6] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[7] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[8] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[9] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[10] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[11] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[12] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[13] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[14] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[15] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[16] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[17] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[18] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[19] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[20] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[21] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[22] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[23] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[24] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[25] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[26] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[27] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[28] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[29] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[2] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[30] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[31] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[3] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[4] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[5] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[6] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[7] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[8] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[9] ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._67_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._69_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._74_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.lzoc_inst._88_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._00_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._00_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._00_[2] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._04_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._04_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._04_[2] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._04_[3] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._10_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._10_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._11_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._14_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._17_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._18_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._22_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._25_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._25_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._25_[2] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._25_[3] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._26_[0] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._26_[1] ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._27_ ;
 wire \sa_inst.cols_l2a:3.l2a_i.rshift._28_[0] ;
 wire \sa_inst.sak._00_[0] ;
 wire \sa_inst.sak._00_[10] ;
 wire \sa_inst.sak._00_[11] ;
 wire \sa_inst.sak._00_[1] ;
 wire \sa_inst.sak._00_[2] ;
 wire \sa_inst.sak._00_[3] ;
 wire \sa_inst.sak._00_[4] ;
 wire \sa_inst.sak._00_[5] ;
 wire \sa_inst.sak._00_[6] ;
 wire \sa_inst.sak._00_[7] ;
 wire \sa_inst.sak._00_[8] ;
 wire \sa_inst.sak._00_[9] ;
 wire \sa_inst.sak._01_[0] ;
 wire \sa_inst.sak._01_[10] ;
 wire \sa_inst.sak._01_[11] ;
 wire \sa_inst.sak._01_[12] ;
 wire \sa_inst.sak._01_[13] ;
 wire \sa_inst.sak._01_[14] ;
 wire \sa_inst.sak._01_[15] ;
 wire \sa_inst.sak._01_[16] ;
 wire \sa_inst.sak._01_[17] ;
 wire \sa_inst.sak._01_[18] ;
 wire \sa_inst.sak._01_[19] ;
 wire \sa_inst.sak._01_[1] ;
 wire \sa_inst.sak._01_[20] ;
 wire \sa_inst.sak._01_[21] ;
 wire \sa_inst.sak._01_[22] ;
 wire \sa_inst.sak._01_[23] ;
 wire \sa_inst.sak._01_[24] ;
 wire \sa_inst.sak._01_[25] ;
 wire \sa_inst.sak._01_[26] ;
 wire \sa_inst.sak._01_[27] ;
 wire \sa_inst.sak._01_[28] ;
 wire \sa_inst.sak._01_[29] ;
 wire \sa_inst.sak._01_[2] ;
 wire \sa_inst.sak._01_[30] ;
 wire \sa_inst.sak._01_[31] ;
 wire \sa_inst.sak._01_[32] ;
 wire \sa_inst.sak._01_[3] ;
 wire \sa_inst.sak._01_[4] ;
 wire \sa_inst.sak._01_[5] ;
 wire \sa_inst.sak._01_[6] ;
 wire \sa_inst.sak._01_[7] ;
 wire \sa_inst.sak._01_[8] ;
 wire \sa_inst.sak._01_[9] ;
 wire \sa_inst.sak._03_[0] ;
 wire \sa_inst.sak._03_[10] ;
 wire \sa_inst.sak._03_[11] ;
 wire \sa_inst.sak._03_[1] ;
 wire \sa_inst.sak._03_[2] ;
 wire \sa_inst.sak._03_[3] ;
 wire \sa_inst.sak._03_[4] ;
 wire \sa_inst.sak._03_[5] ;
 wire \sa_inst.sak._03_[6] ;
 wire \sa_inst.sak._03_[7] ;
 wire \sa_inst.sak._03_[8] ;
 wire \sa_inst.sak._03_[9] ;
 wire \sa_inst.sak._04_ ;
 wire \sa_inst.sak._05_ ;
 wire \sa_inst.sak._06_[0] ;
 wire \sa_inst.sak._06_[10] ;
 wire \sa_inst.sak._06_[11] ;
 wire \sa_inst.sak._06_[12] ;
 wire \sa_inst.sak._06_[13] ;
 wire \sa_inst.sak._06_[14] ;
 wire \sa_inst.sak._06_[15] ;
 wire \sa_inst.sak._06_[16] ;
 wire \sa_inst.sak._06_[17] ;
 wire \sa_inst.sak._06_[18] ;
 wire \sa_inst.sak._06_[19] ;
 wire \sa_inst.sak._06_[1] ;
 wire \sa_inst.sak._06_[20] ;
 wire \sa_inst.sak._06_[21] ;
 wire \sa_inst.sak._06_[22] ;
 wire \sa_inst.sak._06_[23] ;
 wire \sa_inst.sak._06_[24] ;
 wire \sa_inst.sak._06_[25] ;
 wire \sa_inst.sak._06_[26] ;
 wire \sa_inst.sak._06_[27] ;
 wire \sa_inst.sak._06_[28] ;
 wire \sa_inst.sak._06_[29] ;
 wire \sa_inst.sak._06_[2] ;
 wire \sa_inst.sak._06_[30] ;
 wire \sa_inst.sak._06_[31] ;
 wire \sa_inst.sak._06_[32] ;
 wire \sa_inst.sak._06_[3] ;
 wire \sa_inst.sak._06_[4] ;
 wire \sa_inst.sak._06_[5] ;
 wire \sa_inst.sak._06_[6] ;
 wire \sa_inst.sak._06_[7] ;
 wire \sa_inst.sak._06_[8] ;
 wire \sa_inst.sak._06_[9] ;
 wire \sa_inst.sak._07_[0] ;
 wire \sa_inst.sak._07_[10] ;
 wire \sa_inst.sak._07_[11] ;
 wire \sa_inst.sak._07_[1] ;
 wire \sa_inst.sak._07_[2] ;
 wire \sa_inst.sak._07_[3] ;
 wire \sa_inst.sak._07_[4] ;
 wire \sa_inst.sak._07_[5] ;
 wire \sa_inst.sak._07_[6] ;
 wire \sa_inst.sak._07_[7] ;
 wire \sa_inst.sak._07_[8] ;
 wire \sa_inst.sak._07_[9] ;
 wire \sa_inst.sak._08_[0] ;
 wire \sa_inst.sak._08_[10] ;
 wire \sa_inst.sak._08_[11] ;
 wire \sa_inst.sak._08_[1] ;
 wire \sa_inst.sak._08_[2] ;
 wire \sa_inst.sak._08_[3] ;
 wire \sa_inst.sak._08_[4] ;
 wire \sa_inst.sak._08_[5] ;
 wire \sa_inst.sak._08_[6] ;
 wire \sa_inst.sak._08_[7] ;
 wire \sa_inst.sak._08_[8] ;
 wire \sa_inst.sak._08_[9] ;
 wire \sa_inst.sak._09_ ;
 wire \sa_inst.sak._10_ ;
 wire \sa_inst.sak._12_[0] ;
 wire \sa_inst.sak._12_[10] ;
 wire \sa_inst.sak._12_[11] ;
 wire \sa_inst.sak._12_[12] ;
 wire \sa_inst.sak._12_[13] ;
 wire \sa_inst.sak._12_[14] ;
 wire \sa_inst.sak._12_[15] ;
 wire \sa_inst.sak._12_[16] ;
 wire \sa_inst.sak._12_[17] ;
 wire \sa_inst.sak._12_[18] ;
 wire \sa_inst.sak._12_[19] ;
 wire \sa_inst.sak._12_[1] ;
 wire \sa_inst.sak._12_[20] ;
 wire \sa_inst.sak._12_[21] ;
 wire \sa_inst.sak._12_[22] ;
 wire \sa_inst.sak._12_[23] ;
 wire \sa_inst.sak._12_[24] ;
 wire \sa_inst.sak._12_[25] ;
 wire \sa_inst.sak._12_[26] ;
 wire \sa_inst.sak._12_[27] ;
 wire \sa_inst.sak._12_[28] ;
 wire \sa_inst.sak._12_[29] ;
 wire \sa_inst.sak._12_[2] ;
 wire \sa_inst.sak._12_[30] ;
 wire \sa_inst.sak._12_[31] ;
 wire \sa_inst.sak._12_[32] ;
 wire \sa_inst.sak._12_[3] ;
 wire \sa_inst.sak._12_[4] ;
 wire \sa_inst.sak._12_[5] ;
 wire \sa_inst.sak._12_[6] ;
 wire \sa_inst.sak._12_[7] ;
 wire \sa_inst.sak._12_[8] ;
 wire \sa_inst.sak._12_[9] ;
 wire \sa_inst.sak._13_[0] ;
 wire \sa_inst.sak._13_[10] ;
 wire \sa_inst.sak._13_[11] ;
 wire \sa_inst.sak._13_[1] ;
 wire \sa_inst.sak._13_[2] ;
 wire \sa_inst.sak._13_[3] ;
 wire \sa_inst.sak._13_[4] ;
 wire \sa_inst.sak._13_[5] ;
 wire \sa_inst.sak._13_[6] ;
 wire \sa_inst.sak._13_[7] ;
 wire \sa_inst.sak._13_[8] ;
 wire \sa_inst.sak._13_[9] ;
 wire \sa_inst.sak._17_[0] ;
 wire \sa_inst.sak._17_[10] ;
 wire \sa_inst.sak._17_[11] ;
 wire \sa_inst.sak._17_[12] ;
 wire \sa_inst.sak._17_[13] ;
 wire \sa_inst.sak._17_[14] ;
 wire \sa_inst.sak._17_[15] ;
 wire \sa_inst.sak._17_[16] ;
 wire \sa_inst.sak._17_[17] ;
 wire \sa_inst.sak._17_[18] ;
 wire \sa_inst.sak._17_[19] ;
 wire \sa_inst.sak._17_[1] ;
 wire \sa_inst.sak._17_[20] ;
 wire \sa_inst.sak._17_[21] ;
 wire \sa_inst.sak._17_[22] ;
 wire \sa_inst.sak._17_[23] ;
 wire \sa_inst.sak._17_[24] ;
 wire \sa_inst.sak._17_[25] ;
 wire \sa_inst.sak._17_[26] ;
 wire \sa_inst.sak._17_[27] ;
 wire \sa_inst.sak._17_[28] ;
 wire \sa_inst.sak._17_[29] ;
 wire \sa_inst.sak._17_[2] ;
 wire \sa_inst.sak._17_[30] ;
 wire \sa_inst.sak._17_[31] ;
 wire \sa_inst.sak._17_[32] ;
 wire \sa_inst.sak._17_[3] ;
 wire \sa_inst.sak._17_[4] ;
 wire \sa_inst.sak._17_[5] ;
 wire \sa_inst.sak._17_[6] ;
 wire \sa_inst.sak._17_[7] ;
 wire \sa_inst.sak._17_[8] ;
 wire \sa_inst.sak._17_[9] ;
 wire \sa_inst.sak._19_[0] ;
 wire \sa_inst.sak._19_[11] ;
 wire \sa_inst.sak._19_[1] ;
 wire \sa_inst.sak._19_[2] ;
 wire \sa_inst.sak._19_[3] ;
 wire \sa_inst.sak._19_[4] ;
 wire \sa_inst.sak._19_[5] ;
 wire \sa_inst.sak._19_[6] ;
 wire \sa_inst.sak._19_[7] ;
 wire \sa_inst.sak._19_[8] ;
 wire \sa_inst.sak._19_[9] ;
 wire \sa_inst.sak._20_ ;
 wire \sa_inst.sak._21_ ;
 wire \sa_inst.sak._22_ ;
 wire \sa_inst.sak._23_[0] ;
 wire \sa_inst.sak._23_[10] ;
 wire \sa_inst.sak._23_[11] ;
 wire \sa_inst.sak._23_[12] ;
 wire \sa_inst.sak._23_[13] ;
 wire \sa_inst.sak._23_[14] ;
 wire \sa_inst.sak._23_[15] ;
 wire \sa_inst.sak._23_[16] ;
 wire \sa_inst.sak._23_[17] ;
 wire \sa_inst.sak._23_[18] ;
 wire \sa_inst.sak._23_[19] ;
 wire \sa_inst.sak._23_[1] ;
 wire \sa_inst.sak._23_[20] ;
 wire \sa_inst.sak._23_[21] ;
 wire \sa_inst.sak._23_[22] ;
 wire \sa_inst.sak._23_[23] ;
 wire \sa_inst.sak._23_[24] ;
 wire \sa_inst.sak._23_[25] ;
 wire \sa_inst.sak._23_[26] ;
 wire \sa_inst.sak._23_[27] ;
 wire \sa_inst.sak._23_[28] ;
 wire \sa_inst.sak._23_[29] ;
 wire \sa_inst.sak._23_[2] ;
 wire \sa_inst.sak._23_[30] ;
 wire \sa_inst.sak._23_[31] ;
 wire \sa_inst.sak._23_[32] ;
 wire \sa_inst.sak._23_[3] ;
 wire \sa_inst.sak._23_[4] ;
 wire \sa_inst.sak._23_[5] ;
 wire \sa_inst.sak._23_[6] ;
 wire \sa_inst.sak._23_[7] ;
 wire \sa_inst.sak._23_[8] ;
 wire \sa_inst.sak._23_[9] ;
 wire \sa_inst.sak._33_ ;
 wire \sa_inst.sak._40_[0] ;
 wire \sa_inst.sak._40_[10] ;
 wire \sa_inst.sak._40_[11] ;
 wire \sa_inst.sak._40_[12] ;
 wire \sa_inst.sak._40_[13] ;
 wire \sa_inst.sak._40_[14] ;
 wire \sa_inst.sak._40_[15] ;
 wire \sa_inst.sak._40_[16] ;
 wire \sa_inst.sak._40_[17] ;
 wire \sa_inst.sak._40_[18] ;
 wire \sa_inst.sak._40_[19] ;
 wire \sa_inst.sak._40_[1] ;
 wire \sa_inst.sak._40_[20] ;
 wire \sa_inst.sak._40_[21] ;
 wire \sa_inst.sak._40_[22] ;
 wire \sa_inst.sak._40_[23] ;
 wire \sa_inst.sak._40_[24] ;
 wire \sa_inst.sak._40_[25] ;
 wire \sa_inst.sak._40_[26] ;
 wire \sa_inst.sak._40_[27] ;
 wire \sa_inst.sak._40_[28] ;
 wire \sa_inst.sak._40_[29] ;
 wire \sa_inst.sak._40_[2] ;
 wire \sa_inst.sak._40_[30] ;
 wire \sa_inst.sak._40_[31] ;
 wire \sa_inst.sak._40_[32] ;
 wire \sa_inst.sak._40_[3] ;
 wire \sa_inst.sak._40_[4] ;
 wire \sa_inst.sak._40_[5] ;
 wire \sa_inst.sak._40_[6] ;
 wire \sa_inst.sak._40_[7] ;
 wire \sa_inst.sak._40_[8] ;
 wire \sa_inst.sak._40_[9] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[0] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[10] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[11] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[12] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[13] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[14] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[15] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[16] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[17] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[18] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[19] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[1] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[20] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[21] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[22] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[23] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[24] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[25] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[26] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[27] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[28] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[29] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[2] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[30] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[31] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[32] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[3] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[4] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[5] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[6] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[7] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[8] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._00_[9] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._02_ ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[0] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[10] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[11] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[12] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[13] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[14] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[15] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[16] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[17] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[18] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[19] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[1] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[20] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[21] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[22] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[23] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[24] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[25] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[26] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[27] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[28] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[29] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[2] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[30] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[31] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[3] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[4] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[5] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[6] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[7] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[8] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij._10_[9] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._17_ ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._20_ ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[0] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[10] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[11] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[12] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[13] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[14] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[15] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[16] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[17] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[18] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[19] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[1] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[20] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[21] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[22] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[23] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[24] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[25] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[26] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[27] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[28] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[29] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[2] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[30] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[31] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[3] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[4] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[5] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[6] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[7] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[8] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[9] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._25_ ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._26_ ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w10_0 ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w11_0 ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w2_0 ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w3_0 ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w4_0 ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w5_0 ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w6_0 ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w7_0 ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w8_0 ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w9_0 ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ;
 wire \sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[0] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[10] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[11] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[12] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[13] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[14] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[15] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[16] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[17] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[18] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[19] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[1] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[20] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[21] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[22] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[23] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[24] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[25] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[26] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[27] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[28] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[29] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[2] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[30] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[31] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[32] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[3] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[4] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[5] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[6] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[7] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[8] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._00_[9] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._02_ ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[0] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[10] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[11] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[12] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[13] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[14] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[15] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[16] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[17] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[18] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[19] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[1] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[20] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[21] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[22] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[23] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[24] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[25] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[26] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[27] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[28] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[29] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[2] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[30] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[31] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[3] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[4] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[5] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[6] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[7] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[8] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij._10_[9] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._00_ ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._01_ ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._02_ ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._08_[1] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._08_[2] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._08_[3] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._08_[4] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._11_ ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._17_ ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._20_ ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._22_ ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[0] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[10] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[11] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[12] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[13] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[14] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[15] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[16] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[17] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[18] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[19] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[1] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[20] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[21] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[22] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[23] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[24] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[25] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[26] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[27] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[28] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[29] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[2] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[30] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[31] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[3] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[4] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[5] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[6] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[7] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[8] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[9] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._25_ ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._26_ ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[0] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[1] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[2] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[10] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[11] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[12] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[1] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[2] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[3] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[4] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[5] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[6] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[7] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[8] ;
 wire \sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[9] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[0] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[10] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[11] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[12] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[13] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[14] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[15] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[16] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[17] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[18] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[19] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[1] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[20] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[21] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[22] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[23] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[24] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[25] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[26] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[27] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[28] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[29] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[2] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[30] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[31] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[32] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[3] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[4] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[5] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[6] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[7] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[8] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._00_[9] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._02_ ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[0] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[10] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[11] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[12] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[13] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[14] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[15] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[16] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[17] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[18] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[19] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[1] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[20] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[21] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[22] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[23] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[24] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[25] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[26] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[27] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[28] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[29] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[2] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[30] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[31] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[3] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[4] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[5] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[6] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[7] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[8] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij._10_[9] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._00_ ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._01_ ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._02_ ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._08_[1] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._08_[2] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._08_[3] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._08_[4] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._11_ ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._17_ ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._20_ ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._22_ ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[0] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[10] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[11] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[12] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[13] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[14] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[15] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[16] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[17] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[18] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[19] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[1] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[20] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[21] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[22] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[23] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[24] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[25] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[26] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[27] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[28] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[29] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[2] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[30] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[31] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[3] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[4] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[5] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[6] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[7] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[8] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[9] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._25_ ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._26_ ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[0] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[1] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[2] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[10] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[11] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[12] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[1] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[2] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[3] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[4] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[5] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[6] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[7] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[8] ;
 wire \sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[9] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[0] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[10] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[11] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[12] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[13] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[14] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[15] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[16] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[17] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[18] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[19] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[1] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[20] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[21] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[22] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[23] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[24] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[25] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[26] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[27] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[28] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[29] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[2] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[30] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[31] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[32] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[3] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[4] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[5] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[6] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[7] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[8] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._00_[9] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._02_ ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[0] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[10] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[11] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[12] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[13] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[14] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[15] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[16] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[17] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[18] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[19] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[1] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[20] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[21] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[22] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[23] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[24] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[25] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[26] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[27] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[28] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[29] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[2] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[30] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[31] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[3] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[4] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[5] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[6] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[7] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[8] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij._10_[9] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._20_ ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[0] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[10] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[11] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[12] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[13] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[14] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[15] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[16] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[17] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[18] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[19] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[1] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[20] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[21] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[22] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[23] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[24] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[25] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[26] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[27] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[28] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[29] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[2] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[30] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[31] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[3] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[4] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[5] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[6] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[7] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[8] ;
 wire \sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[9] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[0] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[10] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[11] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[12] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[13] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[14] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[15] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[16] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[17] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[18] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[19] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[1] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[20] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[21] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[22] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[23] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[24] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[25] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[26] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[27] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[28] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[29] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[2] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[30] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[31] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[32] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[3] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[4] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[5] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[6] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[7] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[8] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._00_[9] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._02_ ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[0] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[10] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[11] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[12] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[13] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[14] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[15] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[16] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[17] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[18] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[19] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[1] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[20] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[21] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[22] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[23] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[24] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[25] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[26] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[27] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[28] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[29] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[2] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[30] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[31] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[3] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[4] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[5] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[6] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[7] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[8] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij._10_[9] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._20_ ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[0] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[10] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[11] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[12] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[13] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[14] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[15] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[16] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[17] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[18] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[19] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[1] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[20] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[21] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[22] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[23] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[24] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[25] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[26] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[27] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[28] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[29] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[2] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[30] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[31] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[3] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[4] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[5] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[6] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[7] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[8] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[9] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._25_ ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w10_0 ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w11_0 ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w2_0 ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w3_0 ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w4_0 ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w5_0 ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w6_0 ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w7_0 ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w8_0 ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w9_0 ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ;
 wire \sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[0] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[10] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[11] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[12] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[13] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[14] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[15] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[16] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[17] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[18] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[19] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[1] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[20] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[21] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[22] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[23] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[24] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[25] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[26] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[27] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[28] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[29] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[2] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[30] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[31] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[32] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[3] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[4] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[5] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[6] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[7] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[8] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._00_[9] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._02_ ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[0] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[10] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[11] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[12] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[13] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[14] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[15] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[16] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[17] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[18] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[19] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[1] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[20] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[21] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[22] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[23] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[24] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[25] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[26] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[27] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[28] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[29] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[2] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[30] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[31] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[3] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[4] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[5] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[6] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[7] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[8] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij._10_[9] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._00_ ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._01_ ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._02_ ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._08_[1] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._08_[2] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._08_[3] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._08_[4] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._11_ ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._17_ ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._20_ ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._22_ ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[0] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[10] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[11] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[12] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[13] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[14] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[15] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[16] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[17] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[18] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[19] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[1] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[20] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[21] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[22] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[23] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[24] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[25] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[26] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[27] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[28] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[29] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[2] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[30] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[31] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[3] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[4] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[5] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[6] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[7] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[8] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[9] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._25_ ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._26_ ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[0] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[1] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[2] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[10] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[11] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[12] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[1] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[2] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[3] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[4] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[5] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[6] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[7] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[8] ;
 wire \sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[9] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[0] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[10] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[11] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[12] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[13] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[14] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[15] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[16] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[17] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[18] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[19] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[1] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[20] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[21] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[22] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[23] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[24] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[25] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[26] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[27] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[28] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[29] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[2] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[30] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[31] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[32] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[3] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[4] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[5] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[6] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[7] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[8] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._00_[9] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._02_ ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[0] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[10] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[11] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[12] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[13] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[14] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[15] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[16] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[17] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[18] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[19] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[1] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[20] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[21] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[22] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[23] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[24] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[25] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[26] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[27] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[28] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[29] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[2] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[30] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[31] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[3] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[4] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[5] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[6] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[7] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[8] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij._10_[9] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._20_ ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[0] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[10] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[11] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[12] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[13] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[14] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[15] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[16] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[17] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[18] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[19] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[1] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[20] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[21] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[22] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[23] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[24] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[25] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[26] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[27] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[28] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[29] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[2] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[30] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[31] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[3] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[4] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[5] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[6] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[7] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[8] ;
 wire \sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[9] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[0] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[10] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[11] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[12] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[13] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[14] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[15] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[16] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[17] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[18] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[19] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[1] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[20] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[21] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[22] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[23] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[24] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[25] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[26] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[27] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[28] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[29] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[2] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[30] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[31] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[32] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[3] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[4] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[5] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[6] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[7] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[8] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._00_[9] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._02_ ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[0] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[10] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[11] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[12] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[13] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[14] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[15] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[16] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[17] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[18] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[19] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[1] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[20] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[21] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[22] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[23] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[24] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[25] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[26] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[27] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[28] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[29] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[2] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[30] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[31] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[3] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[4] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[5] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[6] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[7] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[8] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij._10_[9] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._20_ ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[0] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[10] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[11] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[12] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[13] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[14] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[15] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[16] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[17] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[18] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[19] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[1] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[20] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[21] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[22] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[23] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[24] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[25] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[26] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[27] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[28] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[29] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[2] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[30] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[31] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[3] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[4] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[5] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[6] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[7] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[8] ;
 wire \sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[9] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[0] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[10] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[11] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[12] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[13] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[14] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[15] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[16] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[17] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[18] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[19] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[1] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[20] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[21] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[22] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[23] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[24] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[25] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[26] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[27] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[28] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[29] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[2] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[30] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[31] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[32] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[3] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[4] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[5] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[6] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[7] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[8] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._00_[9] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._01_ ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._02_ ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[0] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[10] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[11] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[12] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[13] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[14] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[15] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[16] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[17] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[18] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[19] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[1] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[20] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[21] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[22] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[23] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[24] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[25] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[26] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[27] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[28] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[29] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[2] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[30] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[31] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[3] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[4] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[5] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[6] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[7] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[8] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij._10_[9] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._11_ ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._17_ ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._20_ ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._22_ ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[0] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[10] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[11] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[12] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[13] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[14] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[15] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[16] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[17] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[18] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[19] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[1] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[20] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[21] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[22] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[23] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[24] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[25] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[26] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[27] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[28] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[29] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[2] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[30] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[31] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[3] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[4] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[5] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[6] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[7] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[8] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[9] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._25_ ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._26_ ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w10_0 ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w11_0 ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w2_0 ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w3_0 ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w4_0 ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w5_0 ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w6_0 ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w7_0 ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w8_0 ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w9_0 ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[1] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ;
 wire \sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ;
 wire \shift_register[0] ;
 wire \shift_register[10] ;
 wire \shift_register[11] ;
 wire \shift_register[1] ;
 wire \shift_register[2] ;
 wire \shift_register[3] ;
 wire \shift_register[4] ;
 wire \shift_register[5] ;
 wire \shift_register[6] ;
 wire \shift_register[7] ;
 wire \shift_register[8] ;
 wire \shift_register[9] ;

 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_2 _05896_ (.A(\sa_inst.cols_a2s3:1.a2s3_j._23_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst._05_[1] ));
 sky130_fd_sc_hd__clkinv_2 _05897_ (.A(\sa_inst.cols_a2s3:3.a2s3_j._23_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst._07_[1] ));
 sky130_fd_sc_hd__inv_2 _05898_ (.A(\sa_inst.cols_a2s3:2.a2s3_j._23_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst._06_[1] ));
 sky130_fd_sc_hd__or4_1 _05899_ (.A(\sa_inst.cols_l2a:3.l2a_i._00_ ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[16] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[17] ),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00684_));
 sky130_fd_sc_hd__or3_1 _05900_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[29] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[30] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00685_));
 sky130_fd_sc_hd__or4_1 _05901_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[25] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[26] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[27] ),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00686_));
 sky130_fd_sc_hd__or4_1 _05902_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[21] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[22] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[23] ),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00687_));
 sky130_fd_sc_hd__or3_1 _05903_ (.A(_00685_),
    .B(_00686_),
    .C(_00687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00688_));
 sky130_fd_sc_hd__nor4_1 _05904_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[18] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[19] ),
    .C(_00684_),
    .D(_00688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00689_));
 sky130_fd_sc_hd__and4_1 _05905_ (.A(\sa_inst.cols_l2a:3.l2a_i._00_ ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[16] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[17] ),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00690_));
 sky130_fd_sc_hd__and3_1 _05906_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[29] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[30] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00691_));
 sky130_fd_sc_hd__and4_1 _05907_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[25] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[26] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[27] ),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00692_));
 sky130_fd_sc_hd__and4_1 _05908_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[21] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[22] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[23] ),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00693_));
 sky130_fd_sc_hd__and3_1 _05909_ (.A(_00691_),
    .B(_00692_),
    .C(_00693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00694_));
 sky130_fd_sc_hd__and4_1 _05910_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[18] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[19] ),
    .C(_00690_),
    .D(_00694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00695_));
 sky130_fd_sc_hd__nor2_1 _05911_ (.A(_00689_),
    .B(_00695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00696_));
 sky130_fd_sc_hd__clkinv_2 _05912_ (.A(_00696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00697_));
 sky130_fd_sc_hd__clkbuf_2 _05913_ (.A(_00697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00698_));
 sky130_fd_sc_hd__buf_2 _05914_ (.A(_00698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._31_ ));
 sky130_fd_sc_hd__and4_1 _05915_ (.A(\sa_inst._12_[75] ),
    .B(\sa_inst._12_[76] ),
    .C(\sa_inst._12_[77] ),
    .D(\sa_inst._12_[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00699_));
 sky130_fd_sc_hd__and4_1 _05916_ (.A(\sa_inst._12_[79] ),
    .B(\sa_inst._12_[80] ),
    .C(\sa_inst._12_[81] ),
    .D(\sa_inst._12_[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00700_));
 sky130_fd_sc_hd__and4_1 _05917_ (.A(\sa_inst._12_[87] ),
    .B(\sa_inst._12_[88] ),
    .C(\sa_inst._12_[89] ),
    .D(_00700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00701_));
 sky130_fd_sc_hd__or4_1 _05918_ (.A(\sa_inst._12_[75] ),
    .B(\sa_inst._12_[76] ),
    .C(\sa_inst._12_[77] ),
    .D(\sa_inst._12_[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00702_));
 sky130_fd_sc_hd__or4_1 _05919_ (.A(\sa_inst._12_[79] ),
    .B(\sa_inst._12_[80] ),
    .C(\sa_inst._12_[81] ),
    .D(\sa_inst._12_[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00703_));
 sky130_fd_sc_hd__or4_1 _05920_ (.A(\sa_inst._12_[87] ),
    .B(\sa_inst._12_[88] ),
    .C(\sa_inst._12_[89] ),
    .D(_00703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00704_));
 sky130_fd_sc_hd__nor4_1 _05921_ (.A(\sa_inst._12_[97] ),
    .B(\sa_inst._12_[74] ),
    .C(_00702_),
    .D(_00704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00705_));
 sky130_fd_sc_hd__a41o_1 _05922_ (.A1(\sa_inst._12_[97] ),
    .A2(\sa_inst._12_[74] ),
    .A3(_00699_),
    .A4(_00701_),
    .B1(_00705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00706_));
 sky130_fd_sc_hd__and4_1 _05923_ (.A(\sa_inst._12_[69] ),
    .B(\sa_inst._12_[70] ),
    .C(\sa_inst._12_[71] ),
    .D(\sa_inst._12_[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00707_));
 sky130_fd_sc_hd__and4_1 _05924_ (.A(\sa_inst._12_[97] ),
    .B(\sa_inst._12_[66] ),
    .C(\sa_inst._12_[67] ),
    .D(\sa_inst._12_[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00708_));
 sky130_fd_sc_hd__and4_1 _05925_ (.A(\sa_inst._12_[93] ),
    .B(\sa_inst._12_[94] ),
    .C(\sa_inst._12_[95] ),
    .D(\sa_inst._12_[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00709_));
 sky130_fd_sc_hd__and4_1 _05926_ (.A(\sa_inst._12_[85] ),
    .B(\sa_inst._12_[90] ),
    .C(\sa_inst._12_[91] ),
    .D(\sa_inst._12_[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00710_));
 sky130_fd_sc_hd__and4_1 _05927_ (.A(\sa_inst._12_[73] ),
    .B(\sa_inst._12_[82] ),
    .C(\sa_inst._12_[83] ),
    .D(\sa_inst._12_[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00711_));
 sky130_fd_sc_hd__and3_1 _05928_ (.A(_00709_),
    .B(_00710_),
    .C(_00711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00712_));
 sky130_fd_sc_hd__or4_1 _05929_ (.A(\sa_inst._12_[69] ),
    .B(\sa_inst._12_[70] ),
    .C(\sa_inst._12_[71] ),
    .D(\sa_inst._12_[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00713_));
 sky130_fd_sc_hd__or4_1 _05930_ (.A(\sa_inst._12_[97] ),
    .B(\sa_inst._12_[66] ),
    .C(\sa_inst._12_[67] ),
    .D(\sa_inst._12_[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00714_));
 sky130_fd_sc_hd__or4_1 _05931_ (.A(\sa_inst._12_[93] ),
    .B(\sa_inst._12_[94] ),
    .C(\sa_inst._12_[95] ),
    .D(\sa_inst._12_[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00715_));
 sky130_fd_sc_hd__or4_1 _05932_ (.A(\sa_inst._12_[85] ),
    .B(\sa_inst._12_[90] ),
    .C(\sa_inst._12_[91] ),
    .D(\sa_inst._12_[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00716_));
 sky130_fd_sc_hd__or4_1 _05933_ (.A(\sa_inst._12_[73] ),
    .B(\sa_inst._12_[82] ),
    .C(\sa_inst._12_[83] ),
    .D(\sa_inst._12_[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00717_));
 sky130_fd_sc_hd__or3_1 _05934_ (.A(_00715_),
    .B(_00716_),
    .C(_00717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00718_));
 sky130_fd_sc_hd__nor3_1 _05935_ (.A(_00713_),
    .B(_00714_),
    .C(_00718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00719_));
 sky130_fd_sc_hd__a31o_1 _05936_ (.A1(_00707_),
    .A2(_00708_),
    .A3(_00712_),
    .B1(_00719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00720_));
 sky130_fd_sc_hd__nand2_2 _05937_ (.A(_00706_),
    .B(_00720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00721_));
 sky130_fd_sc_hd__clkbuf_2 _05938_ (.A(_00721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00722_));
 sky130_fd_sc_hd__inv_2 _05939_ (.A(_00722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._23_ ));
 sky130_fd_sc_hd__or4_1 _05940_ (.A(\sa_inst.cols_l2a:2.l2a_i._00_ ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[16] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[17] ),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00723_));
 sky130_fd_sc_hd__or3_1 _05941_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[29] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[30] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00724_));
 sky130_fd_sc_hd__or4_1 _05942_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[25] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[26] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[27] ),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00725_));
 sky130_fd_sc_hd__or4_1 _05943_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[21] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[22] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[23] ),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00726_));
 sky130_fd_sc_hd__or3_1 _05944_ (.A(_00724_),
    .B(_00725_),
    .C(_00726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00727_));
 sky130_fd_sc_hd__nor4_1 _05945_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[18] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[19] ),
    .C(_00723_),
    .D(_00727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00728_));
 sky130_fd_sc_hd__and4_1 _05946_ (.A(\sa_inst.cols_l2a:2.l2a_i._00_ ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[16] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[17] ),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00729_));
 sky130_fd_sc_hd__and3_1 _05947_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[29] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[30] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00730_));
 sky130_fd_sc_hd__and4_1 _05948_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[25] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[26] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[27] ),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00731_));
 sky130_fd_sc_hd__and4_1 _05949_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[21] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[22] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[23] ),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00732_));
 sky130_fd_sc_hd__and3_1 _05950_ (.A(_00730_),
    .B(_00731_),
    .C(_00732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00733_));
 sky130_fd_sc_hd__and4_1 _05951_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[18] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[19] ),
    .C(_00729_),
    .D(_00733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00734_));
 sky130_fd_sc_hd__nor2_1 _05952_ (.A(_00728_),
    .B(_00734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00735_));
 sky130_fd_sc_hd__inv_2 _05953_ (.A(_00735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00736_));
 sky130_fd_sc_hd__clkbuf_2 _05954_ (.A(_00736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00737_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05955_ (.A(_00737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00738_));
 sky130_fd_sc_hd__buf_2 _05956_ (.A(_00738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._31_ ));
 sky130_fd_sc_hd__and4_1 _05957_ (.A(\sa_inst._12_[42] ),
    .B(\sa_inst._12_[43] ),
    .C(\sa_inst._12_[44] ),
    .D(\sa_inst._12_[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00739_));
 sky130_fd_sc_hd__and4_1 _05958_ (.A(\sa_inst._12_[46] ),
    .B(\sa_inst._12_[47] ),
    .C(\sa_inst._12_[48] ),
    .D(\sa_inst._12_[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00740_));
 sky130_fd_sc_hd__and4_1 _05959_ (.A(\sa_inst._12_[54] ),
    .B(\sa_inst._12_[55] ),
    .C(\sa_inst._12_[56] ),
    .D(_00740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00741_));
 sky130_fd_sc_hd__or4_1 _05960_ (.A(\sa_inst._12_[42] ),
    .B(\sa_inst._12_[43] ),
    .C(\sa_inst._12_[44] ),
    .D(\sa_inst._12_[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00742_));
 sky130_fd_sc_hd__or4_1 _05961_ (.A(\sa_inst._12_[46] ),
    .B(\sa_inst._12_[47] ),
    .C(\sa_inst._12_[48] ),
    .D(\sa_inst._12_[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00743_));
 sky130_fd_sc_hd__or4_1 _05962_ (.A(\sa_inst._12_[54] ),
    .B(\sa_inst._12_[55] ),
    .C(\sa_inst._12_[56] ),
    .D(_00743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00744_));
 sky130_fd_sc_hd__nor4_1 _05963_ (.A(\sa_inst._12_[64] ),
    .B(\sa_inst._12_[41] ),
    .C(_00742_),
    .D(_00744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00745_));
 sky130_fd_sc_hd__a41o_1 _05964_ (.A1(\sa_inst._12_[64] ),
    .A2(\sa_inst._12_[41] ),
    .A3(_00739_),
    .A4(_00741_),
    .B1(_00745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00746_));
 sky130_fd_sc_hd__and4_1 _05965_ (.A(\sa_inst._12_[36] ),
    .B(\sa_inst._12_[37] ),
    .C(\sa_inst._12_[38] ),
    .D(\sa_inst._12_[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00747_));
 sky130_fd_sc_hd__and4_1 _05966_ (.A(\sa_inst._12_[64] ),
    .B(\sa_inst._12_[33] ),
    .C(\sa_inst._12_[34] ),
    .D(\sa_inst._12_[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00748_));
 sky130_fd_sc_hd__and4_1 _05967_ (.A(\sa_inst._12_[60] ),
    .B(\sa_inst._12_[61] ),
    .C(\sa_inst._12_[62] ),
    .D(\sa_inst._12_[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00749_));
 sky130_fd_sc_hd__and4_1 _05968_ (.A(\sa_inst._12_[52] ),
    .B(\sa_inst._12_[57] ),
    .C(\sa_inst._12_[58] ),
    .D(\sa_inst._12_[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00750_));
 sky130_fd_sc_hd__and4_1 _05969_ (.A(\sa_inst._12_[40] ),
    .B(\sa_inst._12_[49] ),
    .C(\sa_inst._12_[50] ),
    .D(\sa_inst._12_[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00751_));
 sky130_fd_sc_hd__and3_1 _05970_ (.A(_00749_),
    .B(_00750_),
    .C(_00751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00752_));
 sky130_fd_sc_hd__or4_1 _05971_ (.A(\sa_inst._12_[36] ),
    .B(\sa_inst._12_[37] ),
    .C(\sa_inst._12_[38] ),
    .D(\sa_inst._12_[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00753_));
 sky130_fd_sc_hd__or4_1 _05972_ (.A(\sa_inst._12_[64] ),
    .B(\sa_inst._12_[33] ),
    .C(\sa_inst._12_[34] ),
    .D(\sa_inst._12_[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00754_));
 sky130_fd_sc_hd__or4_1 _05973_ (.A(\sa_inst._12_[60] ),
    .B(\sa_inst._12_[61] ),
    .C(\sa_inst._12_[62] ),
    .D(\sa_inst._12_[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00755_));
 sky130_fd_sc_hd__or4_1 _05974_ (.A(\sa_inst._12_[52] ),
    .B(\sa_inst._12_[57] ),
    .C(\sa_inst._12_[58] ),
    .D(\sa_inst._12_[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00756_));
 sky130_fd_sc_hd__or4_1 _05975_ (.A(\sa_inst._12_[40] ),
    .B(\sa_inst._12_[49] ),
    .C(\sa_inst._12_[50] ),
    .D(\sa_inst._12_[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00757_));
 sky130_fd_sc_hd__or3_1 _05976_ (.A(_00755_),
    .B(_00756_),
    .C(_00757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00758_));
 sky130_fd_sc_hd__nor3_1 _05977_ (.A(_00753_),
    .B(_00754_),
    .C(_00758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00759_));
 sky130_fd_sc_hd__a31o_1 _05978_ (.A1(_00747_),
    .A2(_00748_),
    .A3(_00752_),
    .B1(_00759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00760_));
 sky130_fd_sc_hd__nand2_2 _05979_ (.A(_00746_),
    .B(_00760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00761_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05980_ (.A(_00761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00762_));
 sky130_fd_sc_hd__inv_2 _05981_ (.A(_00762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._23_ ));
 sky130_fd_sc_hd__or4_1 _05982_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[17] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[18] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[19] ),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00763_));
 sky130_fd_sc_hd__or3_1 _05983_ (.A(\sa_inst.cols_l2a:1.l2a_i._00_ ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[16] ),
    .C(_00763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00764_));
 sky130_fd_sc_hd__or4_1 _05984_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[25] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[26] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[27] ),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00765_));
 sky130_fd_sc_hd__or4_1 _05985_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[21] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[22] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[23] ),
    .D(_00765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00766_));
 sky130_fd_sc_hd__or4_1 _05986_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[24] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[29] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[30] ),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00767_));
 sky130_fd_sc_hd__nor3_1 _05987_ (.A(_00764_),
    .B(_00766_),
    .C(_00767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00768_));
 sky130_fd_sc_hd__and4_1 _05988_ (.A(\sa_inst.cols_l2a:1.l2a_i._00_ ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[16] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[17] ),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00769_));
 sky130_fd_sc_hd__and3_1 _05989_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[29] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[30] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00770_));
 sky130_fd_sc_hd__and4_1 _05990_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[25] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[26] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[27] ),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00771_));
 sky130_fd_sc_hd__and4_1 _05991_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[21] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[22] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[23] ),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00772_));
 sky130_fd_sc_hd__and3_1 _05992_ (.A(_00770_),
    .B(_00771_),
    .C(_00772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00773_));
 sky130_fd_sc_hd__and4_1 _05993_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[18] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[19] ),
    .C(_00769_),
    .D(_00773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00774_));
 sky130_fd_sc_hd__nor2_1 _05994_ (.A(_00768_),
    .B(_00774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00775_));
 sky130_fd_sc_hd__inv_2 _05995_ (.A(_00775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00776_));
 sky130_fd_sc_hd__clkbuf_2 _05996_ (.A(_00776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00777_));
 sky130_fd_sc_hd__clkbuf_2 _05997_ (.A(_00777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00778_));
 sky130_fd_sc_hd__clkbuf_2 _05998_ (.A(_00778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._31_ ));
 sky130_fd_sc_hd__or4_1 _05999_ (.A(\sa_inst._12_[9] ),
    .B(\sa_inst._12_[10] ),
    .C(\sa_inst._12_[11] ),
    .D(\sa_inst._12_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00779_));
 sky130_fd_sc_hd__or4_1 _06000_ (.A(\sa_inst._12_[13] ),
    .B(\sa_inst._12_[14] ),
    .C(\sa_inst._12_[15] ),
    .D(\sa_inst._12_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00780_));
 sky130_fd_sc_hd__or4_1 _06001_ (.A(\sa_inst._12_[21] ),
    .B(\sa_inst._12_[22] ),
    .C(\sa_inst._12_[23] ),
    .D(_00780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00781_));
 sky130_fd_sc_hd__nor4_2 _06002_ (.A(\sa_inst._12_[31] ),
    .B(\sa_inst._12_[8] ),
    .C(_00779_),
    .D(_00781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00782_));
 sky130_fd_sc_hd__and4_1 _06003_ (.A(\sa_inst._12_[9] ),
    .B(\sa_inst._12_[10] ),
    .C(\sa_inst._12_[11] ),
    .D(\sa_inst._12_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00783_));
 sky130_fd_sc_hd__and4_1 _06004_ (.A(\sa_inst._12_[13] ),
    .B(\sa_inst._12_[14] ),
    .C(\sa_inst._12_[15] ),
    .D(\sa_inst._12_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00784_));
 sky130_fd_sc_hd__and4_1 _06005_ (.A(\sa_inst._12_[21] ),
    .B(\sa_inst._12_[22] ),
    .C(\sa_inst._12_[23] ),
    .D(_00784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00785_));
 sky130_fd_sc_hd__and4_1 _06006_ (.A(\sa_inst._12_[31] ),
    .B(\sa_inst._12_[8] ),
    .C(_00783_),
    .D(_00785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00786_));
 sky130_fd_sc_hd__and4_1 _06007_ (.A(\sa_inst._12_[3] ),
    .B(\sa_inst._12_[4] ),
    .C(\sa_inst._12_[5] ),
    .D(\sa_inst._12_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00787_));
 sky130_fd_sc_hd__and4_1 _06008_ (.A(\sa_inst._12_[31] ),
    .B(\sa_inst._12_[0] ),
    .C(\sa_inst._12_[1] ),
    .D(\sa_inst._12_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00788_));
 sky130_fd_sc_hd__and4_1 _06009_ (.A(\sa_inst._12_[27] ),
    .B(\sa_inst._12_[28] ),
    .C(\sa_inst._12_[29] ),
    .D(\sa_inst._12_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00789_));
 sky130_fd_sc_hd__and4_1 _06010_ (.A(\sa_inst._12_[19] ),
    .B(\sa_inst._12_[24] ),
    .C(\sa_inst._12_[25] ),
    .D(\sa_inst._12_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00790_));
 sky130_fd_sc_hd__and4_1 _06011_ (.A(\sa_inst._12_[7] ),
    .B(\sa_inst._12_[16] ),
    .C(\sa_inst._12_[17] ),
    .D(\sa_inst._12_[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00791_));
 sky130_fd_sc_hd__and3_1 _06012_ (.A(_00789_),
    .B(_00790_),
    .C(_00791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00792_));
 sky130_fd_sc_hd__or4_2 _06013_ (.A(\sa_inst._12_[19] ),
    .B(\sa_inst._12_[24] ),
    .C(\sa_inst._12_[25] ),
    .D(\sa_inst._12_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00793_));
 sky130_fd_sc_hd__or4_1 _06014_ (.A(\sa_inst._12_[27] ),
    .B(\sa_inst._12_[28] ),
    .C(\sa_inst._12_[29] ),
    .D(\sa_inst._12_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00794_));
 sky130_fd_sc_hd__or4_1 _06015_ (.A(\sa_inst._12_[3] ),
    .B(\sa_inst._12_[4] ),
    .C(\sa_inst._12_[5] ),
    .D(\sa_inst._12_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00795_));
 sky130_fd_sc_hd__or4_1 _06016_ (.A(\sa_inst._12_[31] ),
    .B(\sa_inst._12_[0] ),
    .C(\sa_inst._12_[1] ),
    .D(_00795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00796_));
 sky130_fd_sc_hd__or4_1 _06017_ (.A(\sa_inst._12_[16] ),
    .B(\sa_inst._12_[17] ),
    .C(_00794_),
    .D(_00796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00797_));
 sky130_fd_sc_hd__or4_1 _06018_ (.A(\sa_inst._12_[7] ),
    .B(\sa_inst._12_[18] ),
    .C(_00793_),
    .D(_00797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00798_));
 sky130_fd_sc_hd__nor2_1 _06019_ (.A(\sa_inst._12_[2] ),
    .B(_00798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00799_));
 sky130_fd_sc_hd__a31o_1 _06020_ (.A1(_00787_),
    .A2(_00788_),
    .A3(_00792_),
    .B1(_00799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00800_));
 sky130_fd_sc_hd__o21ai_4 _06021_ (.A1(_00782_),
    .A2(_00786_),
    .B1(_00800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00801_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06022_ (.A(_00801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00802_));
 sky130_fd_sc_hd__inv_2 _06023_ (.A(_00802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._23_ ));
 sky130_fd_sc_hd__and4_1 _06024_ (.A(\sa_inst._17_[6] ),
    .B(\sa_inst._17_[2] ),
    .C(\sa_inst._17_[3] ),
    .D(\sa_inst._17_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00803_));
 sky130_fd_sc_hd__nand2_1 _06025_ (.A(\sa_inst._17_[5] ),
    .B(_00803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00804_));
 sky130_fd_sc_hd__or3_1 _06026_ (.A(\sa_inst._17_[6] ),
    .B(\sa_inst._17_[2] ),
    .C(\sa_inst._17_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00805_));
 sky130_fd_sc_hd__or3_1 _06027_ (.A(\sa_inst._17_[3] ),
    .B(\sa_inst._17_[5] ),
    .C(_00805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00806_));
 sky130_fd_sc_hd__nand2_1 _06028_ (.A(_00804_),
    .B(_00806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._11_ ));
 sky130_fd_sc_hd__and4_1 _06029_ (.A(\sa_inst._00_[6] ),
    .B(\sa_inst._00_[2] ),
    .C(\sa_inst._00_[3] ),
    .D(\sa_inst._00_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00807_));
 sky130_fd_sc_hd__nand2_1 _06030_ (.A(\sa_inst._00_[5] ),
    .B(_00807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00808_));
 sky130_fd_sc_hd__or3_1 _06031_ (.A(\sa_inst._00_[6] ),
    .B(\sa_inst._00_[2] ),
    .C(\sa_inst._00_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00809_));
 sky130_fd_sc_hd__or3_1 _06032_ (.A(\sa_inst._00_[3] ),
    .B(\sa_inst._00_[5] ),
    .C(_00809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00810_));
 sky130_fd_sc_hd__nand2_1 _06033_ (.A(_00808_),
    .B(_00810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._11_ ));
 sky130_fd_sc_hd__and2_1 _06034_ (.A(net28),
    .B(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00811_));
 sky130_fd_sc_hd__clkbuf_1 _06035_ (.A(_00811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00812_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06036_ (.A(_00812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00813_));
 sky130_fd_sc_hd__nand2_2 _06037_ (.A(net23),
    .B(_00813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00814_));
 sky130_fd_sc_hd__inv_2 _06038_ (.A(_00814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.arith_in_col_0[6] ));
 sky130_fd_sc_hd__o21a_1 _06039_ (.A1(net17),
    .A2(net23),
    .B1(_00811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00815_));
 sky130_fd_sc_hd__o31a_1 _06040_ (.A1(net20),
    .A2(net21),
    .A3(net22),
    .B1(_00812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00816_));
 sky130_fd_sc_hd__nor2_1 _06041_ (.A(_00815_),
    .B(_00816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00817_));
 sky130_fd_sc_hd__and3_1 _06042_ (.A(net17),
    .B(net21),
    .C(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00818_));
 sky130_fd_sc_hd__and4_1 _06043_ (.A(net23),
    .B(net20),
    .C(_00812_),
    .D(_00818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00819_));
 sky130_fd_sc_hd__nor2_1 _06044_ (.A(_00817_),
    .B(_00819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00820_));
 sky130_fd_sc_hd__inv_2 _06045_ (.A(_00820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._11_ ));
 sky130_fd_sc_hd__mux2_1 _06046_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[3] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[1] ),
    .S(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_1 _06047_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[2] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[0] ),
    .S(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00822_));
 sky130_fd_sc_hd__mux2_1 _06048_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[9] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[7] ),
    .S(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00823_));
 sky130_fd_sc_hd__xnor2_2 _06049_ (.A(\sa_inst.cols_l2a:3.l2a_i._22_ ),
    .B(_00823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00824_));
 sky130_fd_sc_hd__mux2_1 _06050_ (.A0(_00821_),
    .A1(_00822_),
    .S(_00824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00825_));
 sky130_fd_sc_hd__clkbuf_1 _06051_ (.A(_00825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._29_[0] ));
 sky130_fd_sc_hd__mux2_1 _06052_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[4] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[2] ),
    .S(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _06053_ (.A0(_00826_),
    .A1(_00821_),
    .S(_00824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00827_));
 sky130_fd_sc_hd__clkbuf_1 _06054_ (.A(_00827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._29_[1] ));
 sky130_fd_sc_hd__clkbuf_2 _06055_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _06056_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[5] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[3] ),
    .S(_00828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00829_));
 sky130_fd_sc_hd__clkbuf_2 _06057_ (.A(_00824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _06058_ (.A0(_00829_),
    .A1(_00826_),
    .S(_00830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00831_));
 sky130_fd_sc_hd__clkbuf_1 _06059_ (.A(_00831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._29_[2] ));
 sky130_fd_sc_hd__mux2_1 _06060_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[6] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[4] ),
    .S(_00828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00832_));
 sky130_fd_sc_hd__mux2_1 _06061_ (.A0(_00832_),
    .A1(_00829_),
    .S(_00830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00833_));
 sky130_fd_sc_hd__clkbuf_1 _06062_ (.A(_00833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._29_[3] ));
 sky130_fd_sc_hd__mux2_1 _06063_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[7] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[5] ),
    .S(_00828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _06064_ (.A0(_00834_),
    .A1(_00832_),
    .S(_00830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00835_));
 sky130_fd_sc_hd__clkbuf_1 _06065_ (.A(_00835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._29_[4] ));
 sky130_fd_sc_hd__mux2_1 _06066_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[8] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[6] ),
    .S(_00828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _06067_ (.A0(_00836_),
    .A1(_00834_),
    .S(_00830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00837_));
 sky130_fd_sc_hd__clkbuf_1 _06068_ (.A(_00837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._29_[5] ));
 sky130_fd_sc_hd__mux2_1 _06069_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[30] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[22] ),
    .S(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _06070_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[27] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[19] ),
    .S(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _06071_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[28] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[20] ),
    .S(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00840_));
 sky130_fd_sc_hd__clkbuf_2 _06072_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _06073_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[29] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[21] ),
    .S(_00841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00842_));
 sky130_fd_sc_hd__and4_1 _06074_ (.A(\sa_inst.cols_l2a:3.l2a_i._11_ ),
    .B(_00839_),
    .C(_00840_),
    .D(_00842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00843_));
 sky130_fd_sc_hd__or4_1 _06075_ (.A(\sa_inst.cols_l2a:3.l2a_i._11_ ),
    .B(_00838_),
    .C(_00839_),
    .D(_00840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00844_));
 sky130_fd_sc_hd__nor2_1 _06076_ (.A(_00842_),
    .B(_00844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00845_));
 sky130_fd_sc_hd__a21oi_1 _06077_ (.A1(_00838_),
    .A2(_00843_),
    .B1(_00845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00846_));
 sky130_fd_sc_hd__clkbuf_2 _06078_ (.A(_00846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00847_));
 sky130_fd_sc_hd__inv_2 _06079_ (.A(_00847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._56_ ));
 sky130_fd_sc_hd__clkbuf_2 _06080_ (.A(_00841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _06081_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[17] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[9] ),
    .S(_00848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _06082_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[21] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[13] ),
    .S(_00841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _06083_ (.A0(_00849_),
    .A1(_00850_),
    .S(_00847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00851_));
 sky130_fd_sc_hd__clkbuf_1 _06084_ (.A(_00851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[0] ));
 sky130_fd_sc_hd__mux2_1 _06085_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[18] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[10] ),
    .S(_00848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _06086_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[22] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[14] ),
    .S(_00841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _06087_ (.A0(_00852_),
    .A1(_00853_),
    .S(_00847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00854_));
 sky130_fd_sc_hd__clkbuf_1 _06088_ (.A(_00854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[1] ));
 sky130_fd_sc_hd__or2_1 _06089_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[0] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00855_));
 sky130_fd_sc_hd__clkbuf_1 _06090_ (.A(_00855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._74_ ));
 sky130_fd_sc_hd__clkbuf_1 _06091_ (.A(_00696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00856_));
 sky130_fd_sc_hd__and2_1 _06092_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[9] ),
    .B(_00856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00857_));
 sky130_fd_sc_hd__clkbuf_1 _06093_ (.A(_00857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[8] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06094_ (.A(_00856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00858_));
 sky130_fd_sc_hd__and2_1 _06095_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[10] ),
    .B(_00858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00859_));
 sky130_fd_sc_hd__clkbuf_1 _06096_ (.A(_00859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[9] ));
 sky130_fd_sc_hd__and2_1 _06097_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[11] ),
    .B(_00858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00860_));
 sky130_fd_sc_hd__clkbuf_1 _06098_ (.A(_00860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[10] ));
 sky130_fd_sc_hd__and2_1 _06099_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[12] ),
    .B(_00858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00861_));
 sky130_fd_sc_hd__clkbuf_1 _06100_ (.A(_00861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[11] ));
 sky130_fd_sc_hd__and2_1 _06101_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[13] ),
    .B(_00856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00862_));
 sky130_fd_sc_hd__clkbuf_1 _06102_ (.A(_00862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[12] ));
 sky130_fd_sc_hd__and2_1 _06103_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[14] ),
    .B(_00856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00863_));
 sky130_fd_sc_hd__clkbuf_1 _06104_ (.A(_00863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[13] ));
 sky130_fd_sc_hd__and2_1 _06105_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[15] ),
    .B(_00856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00864_));
 sky130_fd_sc_hd__clkbuf_1 _06106_ (.A(_00864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[14] ));
 sky130_fd_sc_hd__mux2_1 _06107_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[16] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._03_ ),
    .S(_00698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00865_));
 sky130_fd_sc_hd__clkbuf_1 _06108_ (.A(_00865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[15] ));
 sky130_fd_sc_hd__or4_1 _06109_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[5] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[6] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[7] ),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00866_));
 sky130_fd_sc_hd__or4_1 _06110_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[1] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[2] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[3] ),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00867_));
 sky130_fd_sc_hd__o21a_1 _06111_ (.A1(_00866_),
    .A2(_00867_),
    .B1(_00858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._50_ ));
 sky130_fd_sc_hd__or4_1 _06112_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[12] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[13] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[14] ),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._50_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00868_));
 sky130_fd_sc_hd__or4_1 _06113_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[8] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[9] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[10] ),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00869_));
 sky130_fd_sc_hd__or3_1 _06114_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[15] ),
    .B(_00868_),
    .C(_00869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00870_));
 sky130_fd_sc_hd__clkbuf_1 _06115_ (.A(_00870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._48_ ));
 sky130_fd_sc_hd__mux2_1 _06116_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[3] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[1] ),
    .S(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _06117_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[2] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[0] ),
    .S(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _06118_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[9] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[7] ),
    .S(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00873_));
 sky130_fd_sc_hd__xnor2_2 _06119_ (.A(\sa_inst.cols_l2a:2.l2a_i._22_ ),
    .B(_00873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00874_));
 sky130_fd_sc_hd__mux2_1 _06120_ (.A0(_00871_),
    .A1(_00872_),
    .S(_00874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00875_));
 sky130_fd_sc_hd__clkbuf_1 _06121_ (.A(_00875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._29_[0] ));
 sky130_fd_sc_hd__mux2_1 _06122_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[4] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[2] ),
    .S(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _06123_ (.A0(_00876_),
    .A1(_00871_),
    .S(_00874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00877_));
 sky130_fd_sc_hd__clkbuf_1 _06124_ (.A(_00877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._29_[1] ));
 sky130_fd_sc_hd__clkbuf_2 _06125_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _06126_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[5] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[3] ),
    .S(_00878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00879_));
 sky130_fd_sc_hd__clkbuf_2 _06127_ (.A(_00874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_1 _06128_ (.A0(_00879_),
    .A1(_00876_),
    .S(_00880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00881_));
 sky130_fd_sc_hd__clkbuf_1 _06129_ (.A(_00881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._29_[2] ));
 sky130_fd_sc_hd__mux2_1 _06130_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[6] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[4] ),
    .S(_00878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00882_));
 sky130_fd_sc_hd__mux2_1 _06131_ (.A0(_00882_),
    .A1(_00879_),
    .S(_00880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00883_));
 sky130_fd_sc_hd__clkbuf_1 _06132_ (.A(_00883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._29_[3] ));
 sky130_fd_sc_hd__mux2_1 _06133_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[7] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[5] ),
    .S(_00878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _06134_ (.A0(_00884_),
    .A1(_00882_),
    .S(_00880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00885_));
 sky130_fd_sc_hd__clkbuf_1 _06135_ (.A(_00885_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._29_[4] ));
 sky130_fd_sc_hd__mux2_1 _06136_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[8] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[6] ),
    .S(_00878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _06137_ (.A0(_00886_),
    .A1(_00884_),
    .S(_00880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00887_));
 sky130_fd_sc_hd__clkbuf_1 _06138_ (.A(_00887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._29_[5] ));
 sky130_fd_sc_hd__mux2_1 _06139_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[30] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[22] ),
    .S(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _06140_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[27] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[19] ),
    .S(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _06141_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[28] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[20] ),
    .S(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00890_));
 sky130_fd_sc_hd__clkbuf_2 _06142_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_1 _06143_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[29] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[21] ),
    .S(_00891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00892_));
 sky130_fd_sc_hd__and4_1 _06144_ (.A(\sa_inst.cols_l2a:2.l2a_i._11_ ),
    .B(_00889_),
    .C(_00890_),
    .D(_00892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00893_));
 sky130_fd_sc_hd__or4_1 _06145_ (.A(\sa_inst.cols_l2a:2.l2a_i._11_ ),
    .B(_00888_),
    .C(_00889_),
    .D(_00890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00894_));
 sky130_fd_sc_hd__nor2_1 _06146_ (.A(_00892_),
    .B(_00894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00895_));
 sky130_fd_sc_hd__a21oi_1 _06147_ (.A1(_00888_),
    .A2(_00893_),
    .B1(_00895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00896_));
 sky130_fd_sc_hd__clkbuf_2 _06148_ (.A(_00896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00897_));
 sky130_fd_sc_hd__inv_2 _06149_ (.A(_00897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._56_ ));
 sky130_fd_sc_hd__clkbuf_2 _06150_ (.A(_00891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _06151_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[17] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[9] ),
    .S(_00898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _06152_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[21] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[13] ),
    .S(_00891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _06153_ (.A0(_00899_),
    .A1(_00900_),
    .S(_00897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00901_));
 sky130_fd_sc_hd__clkbuf_1 _06154_ (.A(_00901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[0] ));
 sky130_fd_sc_hd__mux2_1 _06155_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[18] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[10] ),
    .S(_00898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_1 _06156_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[22] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[14] ),
    .S(_00891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _06157_ (.A0(_00902_),
    .A1(_00903_),
    .S(_00897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00904_));
 sky130_fd_sc_hd__clkbuf_1 _06158_ (.A(_00904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[1] ));
 sky130_fd_sc_hd__or2_1 _06159_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[0] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00905_));
 sky130_fd_sc_hd__clkbuf_1 _06160_ (.A(_00905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._74_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06161_ (.A(_00735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00906_));
 sky130_fd_sc_hd__and2_1 _06162_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[9] ),
    .B(_00906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00907_));
 sky130_fd_sc_hd__clkbuf_1 _06163_ (.A(_00907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[8] ));
 sky130_fd_sc_hd__clkbuf_1 _06164_ (.A(_00906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00908_));
 sky130_fd_sc_hd__and2_1 _06165_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[10] ),
    .B(_00908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00909_));
 sky130_fd_sc_hd__clkbuf_1 _06166_ (.A(_00909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[9] ));
 sky130_fd_sc_hd__and2_1 _06167_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[11] ),
    .B(_00908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00910_));
 sky130_fd_sc_hd__clkbuf_1 _06168_ (.A(_00910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[10] ));
 sky130_fd_sc_hd__and2_1 _06169_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[12] ),
    .B(_00908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00911_));
 sky130_fd_sc_hd__clkbuf_1 _06170_ (.A(_00911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[11] ));
 sky130_fd_sc_hd__and2_1 _06171_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[13] ),
    .B(_00906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00912_));
 sky130_fd_sc_hd__clkbuf_1 _06172_ (.A(_00912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[12] ));
 sky130_fd_sc_hd__and2_1 _06173_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[14] ),
    .B(_00906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00913_));
 sky130_fd_sc_hd__clkbuf_1 _06174_ (.A(_00913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[13] ));
 sky130_fd_sc_hd__and2_1 _06175_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[15] ),
    .B(_00906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00914_));
 sky130_fd_sc_hd__clkbuf_1 _06176_ (.A(_00914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[14] ));
 sky130_fd_sc_hd__mux2_1 _06177_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[16] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._03_ ),
    .S(_00737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00915_));
 sky130_fd_sc_hd__clkbuf_1 _06178_ (.A(_00915_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[15] ));
 sky130_fd_sc_hd__or4_1 _06179_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[5] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[6] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[7] ),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00916_));
 sky130_fd_sc_hd__or4_1 _06180_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[1] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[2] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[3] ),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00917_));
 sky130_fd_sc_hd__o21a_1 _06181_ (.A1(_00916_),
    .A2(_00917_),
    .B1(_00908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._50_ ));
 sky130_fd_sc_hd__or4_1 _06182_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[12] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[13] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[14] ),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._50_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00918_));
 sky130_fd_sc_hd__or4_1 _06183_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[8] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[9] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[10] ),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00919_));
 sky130_fd_sc_hd__or3_1 _06184_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[15] ),
    .B(_00918_),
    .C(_00919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00920_));
 sky130_fd_sc_hd__clkbuf_1 _06185_ (.A(_00920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._48_ ));
 sky130_fd_sc_hd__mux2_1 _06186_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[3] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[1] ),
    .S(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _06187_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[2] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[0] ),
    .S(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _06188_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[9] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[7] ),
    .S(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00923_));
 sky130_fd_sc_hd__xnor2_1 _06189_ (.A(\sa_inst.cols_l2a:1.l2a_i._22_ ),
    .B(_00923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00924_));
 sky130_fd_sc_hd__mux2_1 _06190_ (.A0(_00921_),
    .A1(_00922_),
    .S(_00924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00925_));
 sky130_fd_sc_hd__clkbuf_1 _06191_ (.A(_00925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._29_[0] ));
 sky130_fd_sc_hd__mux2_1 _06192_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[4] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[2] ),
    .S(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _06193_ (.A0(_00926_),
    .A1(_00921_),
    .S(_00924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00927_));
 sky130_fd_sc_hd__clkbuf_1 _06194_ (.A(_00927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._29_[1] ));
 sky130_fd_sc_hd__clkbuf_2 _06195_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _06196_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[5] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[3] ),
    .S(_00928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00929_));
 sky130_fd_sc_hd__clkbuf_2 _06197_ (.A(_00924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _06198_ (.A0(_00929_),
    .A1(_00926_),
    .S(_00930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00931_));
 sky130_fd_sc_hd__clkbuf_1 _06199_ (.A(_00931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._29_[2] ));
 sky130_fd_sc_hd__mux2_1 _06200_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[6] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[4] ),
    .S(_00928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _06201_ (.A0(_00932_),
    .A1(_00929_),
    .S(_00930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00933_));
 sky130_fd_sc_hd__clkbuf_1 _06202_ (.A(_00933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._29_[3] ));
 sky130_fd_sc_hd__mux2_1 _06203_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[7] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[5] ),
    .S(_00928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_1 _06204_ (.A0(_00934_),
    .A1(_00932_),
    .S(_00930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00935_));
 sky130_fd_sc_hd__clkbuf_1 _06205_ (.A(_00935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._29_[4] ));
 sky130_fd_sc_hd__mux2_1 _06206_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[8] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[6] ),
    .S(_00928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _06207_ (.A0(_00936_),
    .A1(_00934_),
    .S(_00930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00937_));
 sky130_fd_sc_hd__clkbuf_1 _06208_ (.A(_00937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._29_[5] ));
 sky130_fd_sc_hd__mux2_1 _06209_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[30] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[22] ),
    .S(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _06210_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[27] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[19] ),
    .S(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _06211_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[28] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[20] ),
    .S(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00940_));
 sky130_fd_sc_hd__clkbuf_2 _06212_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _06213_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[29] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[21] ),
    .S(_00941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00942_));
 sky130_fd_sc_hd__and4_1 _06214_ (.A(\sa_inst.cols_l2a:1.l2a_i._11_ ),
    .B(_00939_),
    .C(_00940_),
    .D(_00942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00943_));
 sky130_fd_sc_hd__or4_1 _06215_ (.A(\sa_inst.cols_l2a:1.l2a_i._11_ ),
    .B(_00938_),
    .C(_00939_),
    .D(_00940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00944_));
 sky130_fd_sc_hd__nor2_1 _06216_ (.A(_00942_),
    .B(_00944_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00945_));
 sky130_fd_sc_hd__a21oi_1 _06217_ (.A1(_00938_),
    .A2(_00943_),
    .B1(_00945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00946_));
 sky130_fd_sc_hd__clkbuf_2 _06218_ (.A(_00946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00947_));
 sky130_fd_sc_hd__inv_2 _06219_ (.A(_00947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._56_ ));
 sky130_fd_sc_hd__clkbuf_2 _06220_ (.A(_00941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _06221_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[17] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[9] ),
    .S(_00948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _06222_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[21] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[13] ),
    .S(_00941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _06223_ (.A0(_00949_),
    .A1(_00950_),
    .S(_00947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00951_));
 sky130_fd_sc_hd__clkbuf_1 _06224_ (.A(_00951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[0] ));
 sky130_fd_sc_hd__mux2_1 _06225_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[18] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[10] ),
    .S(_00948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _06226_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[22] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[14] ),
    .S(_00941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _06227_ (.A0(_00952_),
    .A1(_00953_),
    .S(_00947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00954_));
 sky130_fd_sc_hd__clkbuf_1 _06228_ (.A(_00954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[1] ));
 sky130_fd_sc_hd__or2_1 _06229_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[0] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00955_));
 sky130_fd_sc_hd__clkbuf_1 _06230_ (.A(_00955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._74_ ));
 sky130_fd_sc_hd__clkbuf_1 _06231_ (.A(_00775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00956_));
 sky130_fd_sc_hd__and2_1 _06232_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[9] ),
    .B(_00956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00957_));
 sky130_fd_sc_hd__clkbuf_1 _06233_ (.A(_00957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[8] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06234_ (.A(_00956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00958_));
 sky130_fd_sc_hd__and2_1 _06235_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[10] ),
    .B(_00958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00959_));
 sky130_fd_sc_hd__clkbuf_1 _06236_ (.A(_00959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[9] ));
 sky130_fd_sc_hd__and2_1 _06237_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[11] ),
    .B(_00958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00960_));
 sky130_fd_sc_hd__clkbuf_1 _06238_ (.A(_00960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[10] ));
 sky130_fd_sc_hd__and2_1 _06239_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[12] ),
    .B(_00958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00961_));
 sky130_fd_sc_hd__clkbuf_1 _06240_ (.A(_00961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[11] ));
 sky130_fd_sc_hd__and2_1 _06241_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[13] ),
    .B(_00956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00962_));
 sky130_fd_sc_hd__clkbuf_1 _06242_ (.A(_00962_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[12] ));
 sky130_fd_sc_hd__and2_1 _06243_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[14] ),
    .B(_00956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00963_));
 sky130_fd_sc_hd__clkbuf_1 _06244_ (.A(_00963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[13] ));
 sky130_fd_sc_hd__and2_1 _06245_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[15] ),
    .B(_00956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00964_));
 sky130_fd_sc_hd__clkbuf_1 _06246_ (.A(_00964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[14] ));
 sky130_fd_sc_hd__mux2_1 _06247_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[16] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._03_ ),
    .S(_00777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00965_));
 sky130_fd_sc_hd__clkbuf_1 _06248_ (.A(_00965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[15] ));
 sky130_fd_sc_hd__or4_1 _06249_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[5] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[6] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[7] ),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00966_));
 sky130_fd_sc_hd__or4_1 _06250_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[1] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[2] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[3] ),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00967_));
 sky130_fd_sc_hd__o21a_1 _06251_ (.A1(_00966_),
    .A2(_00967_),
    .B1(_00958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._50_ ));
 sky130_fd_sc_hd__or4_1 _06252_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[12] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[13] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[14] ),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._50_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00968_));
 sky130_fd_sc_hd__or4_1 _06253_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[8] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[9] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[10] ),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00969_));
 sky130_fd_sc_hd__or3_1 _06254_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[15] ),
    .B(_00968_),
    .C(_00969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00970_));
 sky130_fd_sc_hd__clkbuf_1 _06255_ (.A(_00970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._48_ ));
 sky130_fd_sc_hd__mux2_1 _06256_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[25] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[17] ),
    .S(_00841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _06257_ (.A0(_00971_),
    .A1(_00842_),
    .S(_00846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00972_));
 sky130_fd_sc_hd__clkbuf_1 _06258_ (.A(_00972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[8] ));
 sky130_fd_sc_hd__nand2_1 _06259_ (.A(_00838_),
    .B(_00843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00973_));
 sky130_fd_sc_hd__mux2_1 _06260_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[26] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[18] ),
    .S(_00848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00974_));
 sky130_fd_sc_hd__a22o_1 _06261_ (.A1(_00838_),
    .A2(_00973_),
    .B1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._56_ ),
    .B2(_00974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[9] ));
 sky130_fd_sc_hd__nor2_1 _06262_ (.A(\sa_inst.cols_l2a:3.l2a_i._11_ ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00975_));
 sky130_fd_sc_hd__and2_1 _06263_ (.A(\sa_inst.cols_l2a:3.l2a_i._11_ ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _06264_ (.A0(_00975_),
    .A1(_00976_),
    .S(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00977_));
 sky130_fd_sc_hd__clkbuf_1 _06265_ (.A(_00977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._69_ ));
 sky130_fd_sc_hd__mux2_1 _06266_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[24] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[8] ),
    .S(_00697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00978_));
 sky130_fd_sc_hd__clkbuf_1 _06267_ (.A(_00978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[23] ));
 sky130_fd_sc_hd__clkbuf_2 _06268_ (.A(_00697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _06269_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[25] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[9] ),
    .S(_00979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00980_));
 sky130_fd_sc_hd__clkbuf_1 _06270_ (.A(_00980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[24] ));
 sky130_fd_sc_hd__mux2_1 _06271_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[26] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[10] ),
    .S(_00697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00981_));
 sky130_fd_sc_hd__clkbuf_1 _06272_ (.A(_00981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[25] ));
 sky130_fd_sc_hd__mux2_1 _06273_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[27] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[11] ),
    .S(_00697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00982_));
 sky130_fd_sc_hd__clkbuf_1 _06274_ (.A(_00982_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[26] ));
 sky130_fd_sc_hd__mux2_1 _06275_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[28] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[12] ),
    .S(_00979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00983_));
 sky130_fd_sc_hd__clkbuf_1 _06276_ (.A(_00983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[27] ));
 sky130_fd_sc_hd__mux2_1 _06277_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[29] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[13] ),
    .S(_00979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00984_));
 sky130_fd_sc_hd__clkbuf_1 _06278_ (.A(_00984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[28] ));
 sky130_fd_sc_hd__mux2_1 _06279_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[30] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[14] ),
    .S(_00979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00985_));
 sky130_fd_sc_hd__clkbuf_1 _06280_ (.A(_00985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[29] ));
 sky130_fd_sc_hd__mux2_1 _06281_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[31] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[15] ),
    .S(_00979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00986_));
 sky130_fd_sc_hd__clkbuf_1 _06282_ (.A(_00986_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[30] ));
 sky130_fd_sc_hd__or4_1 _06283_ (.A(\sa_inst.cols_l2a:3.l2a_i._00_ ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[23] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[25] ),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00987_));
 sky130_fd_sc_hd__or4_1 _06284_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[28] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[29] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[30] ),
    .D(_00987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00988_));
 sky130_fd_sc_hd__and3_1 _06285_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[28] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[29] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00989_));
 sky130_fd_sc_hd__and4_1 _06286_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[24] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[25] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[26] ),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00990_));
 sky130_fd_sc_hd__nand4_1 _06287_ (.A(\sa_inst.cols_l2a:3.l2a_i._00_ ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[23] ),
    .C(_00989_),
    .D(_00990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00991_));
 sky130_fd_sc_hd__o31ai_1 _06288_ (.A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[24] ),
    .A2(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[27] ),
    .A3(_00988_),
    .B1(_00991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._42_ ));
 sky130_fd_sc_hd__mux2_1 _06289_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[25] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[17] ),
    .S(_00891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _06290_ (.A0(_00992_),
    .A1(_00892_),
    .S(_00896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00993_));
 sky130_fd_sc_hd__clkbuf_1 _06291_ (.A(_00993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[8] ));
 sky130_fd_sc_hd__nand2_1 _06292_ (.A(_00888_),
    .B(_00893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00994_));
 sky130_fd_sc_hd__mux2_1 _06293_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[26] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[18] ),
    .S(_00898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00995_));
 sky130_fd_sc_hd__a22o_1 _06294_ (.A1(_00888_),
    .A2(_00994_),
    .B1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._56_ ),
    .B2(_00995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[9] ));
 sky130_fd_sc_hd__nor2_1 _06295_ (.A(\sa_inst.cols_l2a:2.l2a_i._11_ ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00996_));
 sky130_fd_sc_hd__and2_1 _06296_ (.A(\sa_inst.cols_l2a:2.l2a_i._11_ ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _06297_ (.A0(_00996_),
    .A1(_00997_),
    .S(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00998_));
 sky130_fd_sc_hd__clkbuf_1 _06298_ (.A(_00998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._69_ ));
 sky130_fd_sc_hd__mux2_1 _06299_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[24] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[8] ),
    .S(_00736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00999_));
 sky130_fd_sc_hd__clkbuf_1 _06300_ (.A(_00999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[23] ));
 sky130_fd_sc_hd__mux2_1 _06301_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[25] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[9] ),
    .S(_00736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01000_));
 sky130_fd_sc_hd__clkbuf_1 _06302_ (.A(_01000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[24] ));
 sky130_fd_sc_hd__mux2_1 _06303_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[26] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[10] ),
    .S(_00737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01001_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06304_ (.A(_01001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[25] ));
 sky130_fd_sc_hd__mux2_1 _06305_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[27] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[11] ),
    .S(_00738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01002_));
 sky130_fd_sc_hd__clkbuf_1 _06306_ (.A(_01002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[26] ));
 sky130_fd_sc_hd__mux2_1 _06307_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[28] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[12] ),
    .S(_00736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01003_));
 sky130_fd_sc_hd__clkbuf_1 _06308_ (.A(_01003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[27] ));
 sky130_fd_sc_hd__mux2_1 _06309_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[29] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[13] ),
    .S(_00736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01004_));
 sky130_fd_sc_hd__clkbuf_1 _06310_ (.A(_01004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[28] ));
 sky130_fd_sc_hd__mux2_1 _06311_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[30] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[14] ),
    .S(_00737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01005_));
 sky130_fd_sc_hd__clkbuf_1 _06312_ (.A(_01005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[29] ));
 sky130_fd_sc_hd__mux2_1 _06313_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[31] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[15] ),
    .S(_00737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01006_));
 sky130_fd_sc_hd__clkbuf_1 _06314_ (.A(_01006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[30] ));
 sky130_fd_sc_hd__and4_1 _06315_ (.A(\sa_inst.cols_l2a:2.l2a_i._00_ ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[23] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[24] ),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01007_));
 sky130_fd_sc_hd__and4_1 _06316_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[28] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[29] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[30] ),
    .D(_01007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01008_));
 sky130_fd_sc_hd__or4_1 _06317_ (.A(\sa_inst.cols_l2a:2.l2a_i._00_ ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[23] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[24] ),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01009_));
 sky130_fd_sc_hd__or4_1 _06318_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[28] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[29] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[30] ),
    .D(_01009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01010_));
 sky130_fd_sc_hd__nor3_1 _06319_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[25] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[26] ),
    .C(_01010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01011_));
 sky130_fd_sc_hd__a31o_1 _06320_ (.A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[25] ),
    .A2(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[26] ),
    .A3(_01008_),
    .B1(_01011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._42_ ));
 sky130_fd_sc_hd__mux2_1 _06321_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[25] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[17] ),
    .S(_00941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _06322_ (.A0(_01012_),
    .A1(_00942_),
    .S(_00946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01013_));
 sky130_fd_sc_hd__clkbuf_1 _06323_ (.A(_01013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[8] ));
 sky130_fd_sc_hd__nand2_1 _06324_ (.A(_00938_),
    .B(_00943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01014_));
 sky130_fd_sc_hd__mux2_1 _06325_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[26] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[18] ),
    .S(_00948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01015_));
 sky130_fd_sc_hd__a22o_1 _06326_ (.A1(_00938_),
    .A2(_01014_),
    .B1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._56_ ),
    .B2(_01015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[9] ));
 sky130_fd_sc_hd__nor2_1 _06327_ (.A(\sa_inst.cols_l2a:1.l2a_i._11_ ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01016_));
 sky130_fd_sc_hd__and2_1 _06328_ (.A(\sa_inst.cols_l2a:1.l2a_i._11_ ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _06329_ (.A0(_01016_),
    .A1(_01017_),
    .S(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01018_));
 sky130_fd_sc_hd__clkbuf_1 _06330_ (.A(_01018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._69_ ));
 sky130_fd_sc_hd__mux2_1 _06331_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[24] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[8] ),
    .S(_00776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01019_));
 sky130_fd_sc_hd__clkbuf_1 _06332_ (.A(_01019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[23] ));
 sky130_fd_sc_hd__mux2_1 _06333_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[25] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[9] ),
    .S(_00776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01020_));
 sky130_fd_sc_hd__clkbuf_1 _06334_ (.A(_01020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[24] ));
 sky130_fd_sc_hd__mux2_1 _06335_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[26] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[10] ),
    .S(_00777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01021_));
 sky130_fd_sc_hd__clkbuf_1 _06336_ (.A(_01021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[25] ));
 sky130_fd_sc_hd__mux2_1 _06337_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[27] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[11] ),
    .S(_00778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01022_));
 sky130_fd_sc_hd__clkbuf_1 _06338_ (.A(_01022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[26] ));
 sky130_fd_sc_hd__mux2_1 _06339_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[28] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[12] ),
    .S(_00776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01023_));
 sky130_fd_sc_hd__clkbuf_1 _06340_ (.A(_01023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[27] ));
 sky130_fd_sc_hd__mux2_1 _06341_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[29] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[13] ),
    .S(_00776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01024_));
 sky130_fd_sc_hd__clkbuf_1 _06342_ (.A(_01024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[28] ));
 sky130_fd_sc_hd__mux2_1 _06343_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[30] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[14] ),
    .S(_00777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01025_));
 sky130_fd_sc_hd__clkbuf_1 _06344_ (.A(_01025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[29] ));
 sky130_fd_sc_hd__mux2_1 _06345_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[31] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[15] ),
    .S(_00777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01026_));
 sky130_fd_sc_hd__clkbuf_1 _06346_ (.A(_01026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[30] ));
 sky130_fd_sc_hd__and4_1 _06347_ (.A(\sa_inst.cols_l2a:1.l2a_i._00_ ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[23] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[24] ),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01027_));
 sky130_fd_sc_hd__and4_1 _06348_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[28] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[29] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[30] ),
    .D(_01027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01028_));
 sky130_fd_sc_hd__or4_1 _06349_ (.A(\sa_inst.cols_l2a:1.l2a_i._00_ ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[23] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[24] ),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01029_));
 sky130_fd_sc_hd__or4_1 _06350_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[28] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[29] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[30] ),
    .D(_01029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01030_));
 sky130_fd_sc_hd__nor3_1 _06351_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[25] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[26] ),
    .C(_01030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01031_));
 sky130_fd_sc_hd__a31o_1 _06352_ (.A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[25] ),
    .A2(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[26] ),
    .A3(_01028_),
    .B1(_01031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._42_ ));
 sky130_fd_sc_hd__clkbuf_1 _06353_ (.A(_00804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01032_));
 sky130_fd_sc_hd__a22o_1 _06354_ (.A1(\sa_inst._17_[4] ),
    .A2(_01032_),
    .B1(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._11_ ),
    .B2(\sa_inst._17_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._14_[4] ));
 sky130_fd_sc_hd__clkinv_2 _06355_ (.A(\sa_inst._17_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01033_));
 sky130_fd_sc_hd__a2bb2o_1 _06356_ (.A1_N(_01033_),
    .A2_N(_00803_),
    .B1(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._11_ ),
    .B2(\sa_inst._17_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._14_[5] ));
 sky130_fd_sc_hd__nor2_1 _06357_ (.A(\sa_inst._17_[6] ),
    .B(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._14_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01034_));
 sky130_fd_sc_hd__and2_1 _06358_ (.A(\sa_inst._17_[6] ),
    .B(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._14_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _06359_ (.A0(_01034_),
    .A1(_01035_),
    .S(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._14_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01036_));
 sky130_fd_sc_hd__clkbuf_1 _06360_ (.A(_01036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._01_ ));
 sky130_fd_sc_hd__clkbuf_1 _06361_ (.A(_00808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01037_));
 sky130_fd_sc_hd__a22o_1 _06362_ (.A1(\sa_inst._00_[4] ),
    .A2(_01037_),
    .B1(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._11_ ),
    .B2(\sa_inst._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._14_[4] ));
 sky130_fd_sc_hd__clkinv_2 _06363_ (.A(\sa_inst._00_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01038_));
 sky130_fd_sc_hd__a2bb2o_1 _06364_ (.A1_N(_01038_),
    .A2_N(_00807_),
    .B1(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._11_ ),
    .B2(\sa_inst._00_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._14_[5] ));
 sky130_fd_sc_hd__nor2_1 _06365_ (.A(\sa_inst._00_[6] ),
    .B(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._14_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01039_));
 sky130_fd_sc_hd__and2_1 _06366_ (.A(\sa_inst._00_[6] ),
    .B(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._14_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _06367_ (.A0(_01039_),
    .A1(_01040_),
    .S(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._14_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01041_));
 sky130_fd_sc_hd__clkbuf_1 _06368_ (.A(_01041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._01_ ));
 sky130_fd_sc_hd__and3b_1 _06369_ (.A_N(_00819_),
    .B(_00812_),
    .C(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01042_));
 sky130_fd_sc_hd__a31o_1 _06370_ (.A1(net1),
    .A2(_00813_),
    .A3(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._11_ ),
    .B1(_01042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._14_[4] ));
 sky130_fd_sc_hd__and3b_1 _06371_ (.A_N(_00819_),
    .B(_00812_),
    .C(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01043_));
 sky130_fd_sc_hd__a31o_1 _06372_ (.A1(net12),
    .A2(_00813_),
    .A3(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._11_ ),
    .B1(_01043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._14_[5] ));
 sky130_fd_sc_hd__mux2_1 _06373_ (.A0(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._14_[5] ),
    .A1(_00814_),
    .S(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._14_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01044_));
 sky130_fd_sc_hd__o21ba_1 _06374_ (.A1(_00814_),
    .A2(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._14_[5] ),
    .B1_N(_01044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._01_ ));
 sky130_fd_sc_hd__nand2_1 _06375_ (.A(net24),
    .B(_00813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01045_));
 sky130_fd_sc_hd__inv_2 _06376_ (.A(_01045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.arith_in_col_0[7] ));
 sky130_fd_sc_hd__inv_2 _06377_ (.A(\sa_inst.sak._00_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01046_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06378_ (.A(_01046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01047_));
 sky130_fd_sc_hd__inv_2 _06379_ (.A(\sa_inst.sak._00_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01048_));
 sky130_fd_sc_hd__mux4_1 _06380_ (.A0(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .A1(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .A2(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .A3(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .S0(\sa_inst.sak._00_[0] ),
    .S1(\sa_inst.sak._00_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01049_));
 sky130_fd_sc_hd__clkbuf_2 _06381_ (.A(\sa_inst.sak._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _06382_ (.A0(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ),
    .A1(\sa_inst.sak._00_[4] ),
    .S(_01050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01051_));
 sky130_fd_sc_hd__clkbuf_1 _06383_ (.A(\sa_inst.sak._00_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01052_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06384_ (.A(\sa_inst.sak._00_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01053_));
 sky130_fd_sc_hd__and2b_1 _06385_ (.A_N(_01052_),
    .B(_01053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01054_));
 sky130_fd_sc_hd__a22o_1 _06386_ (.A1(_01048_),
    .A2(_01049_),
    .B1(_01051_),
    .B2(_01054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01055_));
 sky130_fd_sc_hd__and2_2 _06387_ (.A(_01047_),
    .B(_01055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01056_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06388_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01057_));
 sky130_fd_sc_hd__clkbuf_4 _06389_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01058_));
 sky130_fd_sc_hd__nand2_1 _06390_ (.A(_01057_),
    .B(_01058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01059_));
 sky130_fd_sc_hd__xnor2_1 _06391_ (.A(_01056_),
    .B(_01059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[0] ));
 sky130_fd_sc_hd__clkbuf_2 _06392_ (.A(_01048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01060_));
 sky130_fd_sc_hd__mux4_2 _06393_ (.A0(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .A1(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .A2(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .A3(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .S0(_01050_),
    .S1(\sa_inst.sak._00_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01061_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06394_ (.A(\sa_inst.sak._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01062_));
 sky130_fd_sc_hd__and2b_1 _06395_ (.A_N(_01062_),
    .B(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01063_));
 sky130_fd_sc_hd__a22o_1 _06396_ (.A1(_01060_),
    .A2(_01061_),
    .B1(_01063_),
    .B2(_01054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01064_));
 sky130_fd_sc_hd__and3_1 _06397_ (.A(_01047_),
    .B(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[1] ),
    .C(_01064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01065_));
 sky130_fd_sc_hd__a21o_1 _06398_ (.A1(_01047_),
    .A2(_01064_),
    .B1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01066_));
 sky130_fd_sc_hd__and2b_1 _06399_ (.A_N(_01065_),
    .B(_01066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01067_));
 sky130_fd_sc_hd__clkinv_2 _06400_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01068_));
 sky130_fd_sc_hd__a31o_1 _06401_ (.A1(_01057_),
    .A2(_01056_),
    .A3(_01067_),
    .B1(_01068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01069_));
 sky130_fd_sc_hd__a21oi_1 _06402_ (.A1(_01057_),
    .A2(_01056_),
    .B1(_01067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01070_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06403_ (.A(_01046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01071_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06404_ (.A(_01071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01072_));
 sky130_fd_sc_hd__and2_1 _06405_ (.A(_01072_),
    .B(_01064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01073_));
 sky130_fd_sc_hd__buf_2 _06406_ (.A(_01068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01074_));
 sky130_fd_sc_hd__a2bb2o_1 _06407_ (.A1_N(_01069_),
    .A2_N(_01070_),
    .B1(_01073_),
    .B2(_01074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[1] ));
 sky130_fd_sc_hd__a31o_1 _06408_ (.A1(_01057_),
    .A2(_01056_),
    .A3(_01066_),
    .B1(_01065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01075_));
 sky130_fd_sc_hd__clkbuf_2 _06409_ (.A(_01053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _06410_ (.A0(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .A1(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .S(_01050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01077_));
 sky130_fd_sc_hd__clkbuf_2 _06411_ (.A(\sa_inst.sak._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01078_));
 sky130_fd_sc_hd__and2_1 _06412_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .B(_01078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01079_));
 sky130_fd_sc_hd__inv_2 _06413_ (.A(\sa_inst.sak._00_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01080_));
 sky130_fd_sc_hd__mux2_2 _06414_ (.A0(_01077_),
    .A1(_01079_),
    .S(_01080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _06415_ (.A0(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .A1(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ),
    .S(_01050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01082_));
 sky130_fd_sc_hd__and3b_1 _06416_ (.A_N(_01062_),
    .B(\sa_inst.sak._00_[4] ),
    .C(_01052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01083_));
 sky130_fd_sc_hd__a211o_1 _06417_ (.A1(_01080_),
    .A2(_01082_),
    .B1(_01083_),
    .C1(_01060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01084_));
 sky130_fd_sc_hd__o211a_1 _06418_ (.A1(_01076_),
    .A2(_01081_),
    .B1(_01084_),
    .C1(_01071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01085_));
 sky130_fd_sc_hd__or2_2 _06419_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[2] ),
    .B(_01085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01086_));
 sky130_fd_sc_hd__nand2_1 _06420_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[2] ),
    .B(_01085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01087_));
 sky130_fd_sc_hd__and3_1 _06421_ (.A(_01075_),
    .B(_01086_),
    .C(_01087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01088_));
 sky130_fd_sc_hd__a21oi_1 _06422_ (.A1(_01086_),
    .A2(_01087_),
    .B1(_01075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01089_));
 sky130_fd_sc_hd__nand2_1 _06423_ (.A(_01074_),
    .B(_01085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01090_));
 sky130_fd_sc_hd__o31ai_1 _06424_ (.A1(_01068_),
    .A2(_01088_),
    .A3(_01089_),
    .B1(_01090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[2] ));
 sky130_fd_sc_hd__mux2_1 _06425_ (.A0(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .A1(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .S(_01050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01091_));
 sky130_fd_sc_hd__and2_1 _06426_ (.A(_01062_),
    .B(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _06427_ (.A0(_01091_),
    .A1(_01092_),
    .S(_01080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _06428_ (.A0(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .A1(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ),
    .S(_01078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01094_));
 sky130_fd_sc_hd__and3_1 _06429_ (.A(_01046_),
    .B(_01054_),
    .C(_01094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01095_));
 sky130_fd_sc_hd__a31o_1 _06430_ (.A1(_01060_),
    .A2(_01047_),
    .A3(_01093_),
    .B1(_01095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01096_));
 sky130_fd_sc_hd__or2_1 _06431_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[3] ),
    .B(_01096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01097_));
 sky130_fd_sc_hd__nand2_1 _06432_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[3] ),
    .B(_01096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01098_));
 sky130_fd_sc_hd__nand2_1 _06433_ (.A(_01097_),
    .B(_01098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01099_));
 sky130_fd_sc_hd__o2111a_1 _06434_ (.A1(_01076_),
    .A2(_01081_),
    .B1(_01084_),
    .C1(_01071_),
    .D1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01100_));
 sky130_fd_sc_hd__a311o_1 _06435_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[0] ),
    .A2(_01056_),
    .A3(_01066_),
    .B1(_01100_),
    .C1(_01065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01101_));
 sky130_fd_sc_hd__nand2_1 _06436_ (.A(_01086_),
    .B(_01101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01102_));
 sky130_fd_sc_hd__xor2_1 _06437_ (.A(_01099_),
    .B(_01102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _06438_ (.A0(_01096_),
    .A1(_01103_),
    .S(_01058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01104_));
 sky130_fd_sc_hd__clkbuf_1 _06439_ (.A(_01104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[3] ));
 sky130_fd_sc_hd__mux2_1 _06440_ (.A0(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .A1(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .S(_01078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01105_));
 sky130_fd_sc_hd__a21o_1 _06441_ (.A1(_01052_),
    .A2(_01105_),
    .B1(_01053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_1 _06442_ (.A0(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .A1(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .S(_01078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01107_));
 sky130_fd_sc_hd__or2b_1 _06443_ (.A(\sa_inst.sak._00_[1] ),
    .B_N(_01053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01108_));
 sky130_fd_sc_hd__nand2_1 _06444_ (.A(_01053_),
    .B(_01052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01109_));
 sky130_fd_sc_hd__o22a_1 _06445_ (.A1(_01107_),
    .A2(_01108_),
    .B1(_01109_),
    .B2(_01051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01110_));
 sky130_fd_sc_hd__and3_1 _06446_ (.A(_01047_),
    .B(_01106_),
    .C(_01110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01111_));
 sky130_fd_sc_hd__and2_1 _06447_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[4] ),
    .B(_01111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01112_));
 sky130_fd_sc_hd__nor2_1 _06448_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[4] ),
    .B(_01111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01113_));
 sky130_fd_sc_hd__or2_1 _06449_ (.A(_01112_),
    .B(_01113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01114_));
 sky130_fd_sc_hd__and2_1 _06450_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[3] ),
    .B(_01096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01115_));
 sky130_fd_sc_hd__a31oi_4 _06451_ (.A1(_01086_),
    .A2(_01097_),
    .A3(_01101_),
    .B1(_01115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01116_));
 sky130_fd_sc_hd__xor2_1 _06452_ (.A(_01114_),
    .B(_01116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _06453_ (.A0(_01111_),
    .A1(_01117_),
    .S(_01058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01118_));
 sky130_fd_sc_hd__clkbuf_1 _06454_ (.A(_01118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[4] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06455_ (.A(_01052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _06456_ (.A0(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .A1(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .S(_01062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01120_));
 sky130_fd_sc_hd__a21o_1 _06457_ (.A1(_01119_),
    .A2(_01120_),
    .B1(_01076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _06458_ (.A0(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .A1(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .S(_01078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01122_));
 sky130_fd_sc_hd__o22a_1 _06459_ (.A1(_01108_),
    .A2(_01122_),
    .B1(_01063_),
    .B2(_01109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01123_));
 sky130_fd_sc_hd__and3_1 _06460_ (.A(_01071_),
    .B(_01121_),
    .C(_01123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01124_));
 sky130_fd_sc_hd__and2_1 _06461_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[5] ),
    .B(_01124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01125_));
 sky130_fd_sc_hd__or2_1 _06462_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[5] ),
    .B(_01124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01126_));
 sky130_fd_sc_hd__or2b_1 _06463_ (.A(_01125_),
    .B_N(_01126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01127_));
 sky130_fd_sc_hd__o21bai_1 _06464_ (.A1(_01114_),
    .A2(_01116_),
    .B1_N(_01112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01128_));
 sky130_fd_sc_hd__xnor2_1 _06465_ (.A(_01127_),
    .B(_01128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01129_));
 sky130_fd_sc_hd__mux2_1 _06466_ (.A0(_01124_),
    .A1(_01129_),
    .S(_01058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01130_));
 sky130_fd_sc_hd__clkbuf_1 _06467_ (.A(_01130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[5] ));
 sky130_fd_sc_hd__o22a_1 _06468_ (.A1(_01108_),
    .A2(_01077_),
    .B1(_01082_),
    .B2(_01109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01131_));
 sky130_fd_sc_hd__clkbuf_4 _06469_ (.A(_01062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01132_));
 sky130_fd_sc_hd__a31o_1 _06470_ (.A1(_01119_),
    .A2(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .A3(_01132_),
    .B1(_01076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01133_));
 sky130_fd_sc_hd__and3_1 _06471_ (.A(_01071_),
    .B(_01131_),
    .C(_01133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01134_));
 sky130_fd_sc_hd__and2_1 _06472_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[6] ),
    .B(_01134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01135_));
 sky130_fd_sc_hd__nor2_1 _06473_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[6] ),
    .B(_01134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01136_));
 sky130_fd_sc_hd__nor2_1 _06474_ (.A(_01135_),
    .B(_01136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01137_));
 sky130_fd_sc_hd__o21ai_1 _06475_ (.A1(_01112_),
    .A2(_01125_),
    .B1(_01126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01138_));
 sky130_fd_sc_hd__o31a_1 _06476_ (.A1(_01114_),
    .A2(_01116_),
    .A3(_01127_),
    .B1(_01138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01139_));
 sky130_fd_sc_hd__xnor2_1 _06477_ (.A(_01137_),
    .B(_01139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01140_));
 sky130_fd_sc_hd__buf_2 _06478_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _06479_ (.A0(_01134_),
    .A1(_01140_),
    .S(_01141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01142_));
 sky130_fd_sc_hd__clkbuf_1 _06480_ (.A(_01142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[6] ));
 sky130_fd_sc_hd__o22a_1 _06481_ (.A1(_01108_),
    .A2(_01091_),
    .B1(_01109_),
    .B2(_01094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01143_));
 sky130_fd_sc_hd__clkbuf_2 _06482_ (.A(_01076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01144_));
 sky130_fd_sc_hd__a31o_1 _06483_ (.A1(_01119_),
    .A2(_01132_),
    .A3(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .B1(_01144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01145_));
 sky130_fd_sc_hd__and3_1 _06484_ (.A(_01072_),
    .B(_01143_),
    .C(_01145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01146_));
 sky130_fd_sc_hd__and2_1 _06485_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[7] ),
    .B(_01146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01147_));
 sky130_fd_sc_hd__nor2_1 _06486_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[7] ),
    .B(_01146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01148_));
 sky130_fd_sc_hd__nor2_1 _06487_ (.A(_01147_),
    .B(_01148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01149_));
 sky130_fd_sc_hd__inv_2 _06488_ (.A(_01137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01150_));
 sky130_fd_sc_hd__o21ba_1 _06489_ (.A1(_01150_),
    .A2(_01139_),
    .B1_N(_01135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01151_));
 sky130_fd_sc_hd__xnor2_1 _06490_ (.A(_01149_),
    .B(_01151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01152_));
 sky130_fd_sc_hd__mux2_1 _06491_ (.A0(_01146_),
    .A1(_01152_),
    .S(_01141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01153_));
 sky130_fd_sc_hd__clkbuf_1 _06492_ (.A(_01153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[7] ));
 sky130_fd_sc_hd__nor2_1 _06493_ (.A(_01135_),
    .B(_01147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01154_));
 sky130_fd_sc_hd__o21a_1 _06494_ (.A1(_01150_),
    .A2(_01139_),
    .B1(_01154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01155_));
 sky130_fd_sc_hd__and3_1 _06495_ (.A(_01144_),
    .B(_01072_),
    .C(_01049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01156_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06496_ (.A(_01156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01157_));
 sky130_fd_sc_hd__xnor2_1 _06497_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[8] ),
    .B(_01157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01158_));
 sky130_fd_sc_hd__o21a_1 _06498_ (.A1(_01148_),
    .A2(_01155_),
    .B1(_01158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01159_));
 sky130_fd_sc_hd__nor3_1 _06499_ (.A(_01148_),
    .B(_01158_),
    .C(_01155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01160_));
 sky130_fd_sc_hd__nand2_1 _06500_ (.A(_01068_),
    .B(_01157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01161_));
 sky130_fd_sc_hd__o31ai_1 _06501_ (.A1(_01068_),
    .A2(_01159_),
    .A3(_01160_),
    .B1(_01161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[8] ));
 sky130_fd_sc_hd__and3_1 _06502_ (.A(_01144_),
    .B(_01072_),
    .C(_01061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01162_));
 sky130_fd_sc_hd__nor2_2 _06503_ (.A(_01060_),
    .B(\sa_inst.sak._00_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01163_));
 sky130_fd_sc_hd__and3_1 _06504_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[9] ),
    .B(_01061_),
    .C(_01163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01164_));
 sky130_fd_sc_hd__nor2_1 _06505_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[9] ),
    .B(_01162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01165_));
 sky130_fd_sc_hd__or2_1 _06506_ (.A(_01164_),
    .B(_01165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01166_));
 sky130_fd_sc_hd__a21oi_1 _06507_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[8] ),
    .A2(_01157_),
    .B1(_01160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01167_));
 sky130_fd_sc_hd__xor2_1 _06508_ (.A(_01166_),
    .B(_01167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _06509_ (.A0(_01162_),
    .A1(_01168_),
    .S(_01141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01169_));
 sky130_fd_sc_hd__clkbuf_1 _06510_ (.A(_01169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[9] ));
 sky130_fd_sc_hd__and2_1 _06511_ (.A(_01081_),
    .B(_01163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01170_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06512_ (.A(_01163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01171_));
 sky130_fd_sc_hd__and3_1 _06513_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[10] ),
    .B(_01081_),
    .C(_01171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01172_));
 sky130_fd_sc_hd__nor2_1 _06514_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[10] ),
    .B(_01170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01173_));
 sky130_fd_sc_hd__or2_1 _06515_ (.A(_01172_),
    .B(_01173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01174_));
 sky130_fd_sc_hd__inv_2 _06516_ (.A(_01165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01175_));
 sky130_fd_sc_hd__a21oi_1 _06517_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[8] ),
    .A2(_01157_),
    .B1(_01164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01176_));
 sky130_fd_sc_hd__o31ai_1 _06518_ (.A1(_01148_),
    .A2(_01158_),
    .A3(_01155_),
    .B1(_01176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01177_));
 sky130_fd_sc_hd__and2_1 _06519_ (.A(_01175_),
    .B(_01177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01178_));
 sky130_fd_sc_hd__xnor2_1 _06520_ (.A(_01174_),
    .B(_01178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01179_));
 sky130_fd_sc_hd__mux2_1 _06521_ (.A0(_01170_),
    .A1(_01179_),
    .S(_01141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01180_));
 sky130_fd_sc_hd__clkbuf_1 _06522_ (.A(_01180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[10] ));
 sky130_fd_sc_hd__and2_1 _06523_ (.A(_01171_),
    .B(_01093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01181_));
 sky130_fd_sc_hd__and3_1 _06524_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[11] ),
    .B(_01171_),
    .C(_01093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01182_));
 sky130_fd_sc_hd__or2_1 _06525_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[11] ),
    .B(_01181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01183_));
 sky130_fd_sc_hd__and2b_1 _06526_ (.A_N(_01182_),
    .B(_01183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01184_));
 sky130_fd_sc_hd__inv_2 _06527_ (.A(_01173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01185_));
 sky130_fd_sc_hd__a21oi_1 _06528_ (.A1(_01185_),
    .A2(_01178_),
    .B1(_01172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01186_));
 sky130_fd_sc_hd__xnor2_1 _06529_ (.A(_01184_),
    .B(_01186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01187_));
 sky130_fd_sc_hd__mux2_1 _06530_ (.A0(_01181_),
    .A1(_01187_),
    .S(_01141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01188_));
 sky130_fd_sc_hd__clkbuf_1 _06531_ (.A(_01188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[11] ));
 sky130_fd_sc_hd__and3_1 _06532_ (.A(_01119_),
    .B(_01105_),
    .C(_01163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01189_));
 sky130_fd_sc_hd__and2_1 _06533_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[12] ),
    .B(_01189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01190_));
 sky130_fd_sc_hd__nor2_1 _06534_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[12] ),
    .B(_01189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01191_));
 sky130_fd_sc_hd__or2_1 _06535_ (.A(_01190_),
    .B(_01191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01192_));
 sky130_fd_sc_hd__a311o_1 _06536_ (.A1(_01175_),
    .A2(_01185_),
    .A3(_01177_),
    .B1(_01182_),
    .C1(_01172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01193_));
 sky130_fd_sc_hd__and2_1 _06537_ (.A(_01183_),
    .B(_01193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01194_));
 sky130_fd_sc_hd__xnor2_1 _06538_ (.A(_01192_),
    .B(_01194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01195_));
 sky130_fd_sc_hd__clkbuf_2 _06539_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _06540_ (.A0(_01189_),
    .A1(_01195_),
    .S(_01196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01197_));
 sky130_fd_sc_hd__clkbuf_1 _06541_ (.A(_01197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[12] ));
 sky130_fd_sc_hd__clkbuf_2 _06542_ (.A(_01196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01198_));
 sky130_fd_sc_hd__buf_2 _06543_ (.A(_01119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01199_));
 sky130_fd_sc_hd__and3_1 _06544_ (.A(_01199_),
    .B(_01120_),
    .C(_01171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01200_));
 sky130_fd_sc_hd__and2_1 _06545_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[13] ),
    .B(_01200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01201_));
 sky130_fd_sc_hd__nor2_1 _06546_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[13] ),
    .B(_01200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01202_));
 sky130_fd_sc_hd__nor2_1 _06547_ (.A(_01201_),
    .B(_01202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01203_));
 sky130_fd_sc_hd__inv_2 _06548_ (.A(_01192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01204_));
 sky130_fd_sc_hd__a31o_1 _06549_ (.A1(_01183_),
    .A2(_01204_),
    .A3(_01193_),
    .B1(_01190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01205_));
 sky130_fd_sc_hd__xnor2_1 _06550_ (.A(_01203_),
    .B(_01205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01206_));
 sky130_fd_sc_hd__clkbuf_2 _06551_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01207_));
 sky130_fd_sc_hd__nor2_1 _06552_ (.A(_01207_),
    .B(_01200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01208_));
 sky130_fd_sc_hd__a21oi_1 _06553_ (.A1(_01198_),
    .A2(_01206_),
    .B1(_01208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[13] ));
 sky130_fd_sc_hd__and3_1 _06554_ (.A(_01199_),
    .B(_01079_),
    .C(_01163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01209_));
 sky130_fd_sc_hd__and2_1 _06555_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[14] ),
    .B(_01209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01210_));
 sky130_fd_sc_hd__nor2_1 _06556_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[14] ),
    .B(_01209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01211_));
 sky130_fd_sc_hd__or2_1 _06557_ (.A(_01210_),
    .B(_01211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01212_));
 sky130_fd_sc_hd__o21ba_1 _06558_ (.A1(_01190_),
    .A2(_01201_),
    .B1_N(_01202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01213_));
 sky130_fd_sc_hd__a41o_1 _06559_ (.A1(_01183_),
    .A2(_01204_),
    .A3(_01193_),
    .A4(_01203_),
    .B1(_01213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01214_));
 sky130_fd_sc_hd__xnor2_1 _06560_ (.A(_01212_),
    .B(_01214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01215_));
 sky130_fd_sc_hd__mux2_1 _06561_ (.A0(_01209_),
    .A1(_01215_),
    .S(_01196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01216_));
 sky130_fd_sc_hd__clkbuf_1 _06562_ (.A(_01216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[14] ));
 sky130_fd_sc_hd__and3_1 _06563_ (.A(_01199_),
    .B(_01171_),
    .C(_01092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01217_));
 sky130_fd_sc_hd__and2_1 _06564_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[15] ),
    .B(_01217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01218_));
 sky130_fd_sc_hd__nor2_1 _06565_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[15] ),
    .B(_01217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01219_));
 sky130_fd_sc_hd__nor2_1 _06566_ (.A(_01218_),
    .B(_01219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01220_));
 sky130_fd_sc_hd__inv_2 _06567_ (.A(_01212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01221_));
 sky130_fd_sc_hd__a21oi_1 _06568_ (.A1(_01221_),
    .A2(_01214_),
    .B1(_01210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01222_));
 sky130_fd_sc_hd__xnor2_1 _06569_ (.A(_01220_),
    .B(_01222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01223_));
 sky130_fd_sc_hd__mux2_1 _06570_ (.A0(_01217_),
    .A1(_01223_),
    .S(_01196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01224_));
 sky130_fd_sc_hd__clkbuf_1 _06571_ (.A(_01224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[15] ));
 sky130_fd_sc_hd__o21ba_1 _06572_ (.A1(_01210_),
    .A2(_01218_),
    .B1_N(_01219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01225_));
 sky130_fd_sc_hd__a31o_1 _06573_ (.A1(_01221_),
    .A2(_01214_),
    .A3(_01220_),
    .B1(_01225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01226_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06574_ (.A(_01226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01227_));
 sky130_fd_sc_hd__a21oi_1 _06575_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[16] ),
    .A2(_01227_),
    .B1(_01074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01228_));
 sky130_fd_sc_hd__o21a_1 _06576_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[16] ),
    .A2(_01227_),
    .B1(_01228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[16] ));
 sky130_fd_sc_hd__and2_1 _06577_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[16] ),
    .B(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01229_));
 sky130_fd_sc_hd__a21oi_1 _06578_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[16] ),
    .A2(_01227_),
    .B1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01230_));
 sky130_fd_sc_hd__a211oi_1 _06579_ (.A1(_01227_),
    .A2(_01229_),
    .B1(_01230_),
    .C1(_01074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[17] ));
 sky130_fd_sc_hd__and3_1 _06580_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[18] ),
    .B(_01226_),
    .C(_01229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01231_));
 sky130_fd_sc_hd__a21o_1 _06581_ (.A1(_01227_),
    .A2(_01229_),
    .B1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01232_));
 sky130_fd_sc_hd__and3b_1 _06582_ (.A_N(_01231_),
    .B(_01207_),
    .C(_01232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01233_));
 sky130_fd_sc_hd__clkbuf_1 _06583_ (.A(_01233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[18] ));
 sky130_fd_sc_hd__and4_1 _06584_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[18] ),
    .B(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[19] ),
    .C(_01226_),
    .D(_01229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01234_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06585_ (.A(_01234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01235_));
 sky130_fd_sc_hd__nor2_1 _06586_ (.A(_01074_),
    .B(_01235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01236_));
 sky130_fd_sc_hd__o21a_1 _06587_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[19] ),
    .A2(_01231_),
    .B1(_01236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[19] ));
 sky130_fd_sc_hd__and2_1 _06588_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[20] ),
    .B(_01235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01237_));
 sky130_fd_sc_hd__o21ai_1 _06589_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[20] ),
    .A2(_01235_),
    .B1(_01198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01238_));
 sky130_fd_sc_hd__nor2_1 _06590_ (.A(_01237_),
    .B(_01238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[20] ));
 sky130_fd_sc_hd__and2_1 _06591_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[20] ),
    .B(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01239_));
 sky130_fd_sc_hd__and2_1 _06592_ (.A(_01235_),
    .B(_01239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01240_));
 sky130_fd_sc_hd__inv_2 _06593_ (.A(_01240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01241_));
 sky130_fd_sc_hd__o211a_1 _06594_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[21] ),
    .A2(_01237_),
    .B1(_01241_),
    .C1(_01198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[21] ));
 sky130_fd_sc_hd__and3_1 _06595_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[22] ),
    .B(_01235_),
    .C(_01239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01242_));
 sky130_fd_sc_hd__o21ai_1 _06596_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[22] ),
    .A2(_01240_),
    .B1(_01198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01243_));
 sky130_fd_sc_hd__nor2_1 _06597_ (.A(_01242_),
    .B(_01243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[22] ));
 sky130_fd_sc_hd__and4_1 _06598_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[22] ),
    .B(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[23] ),
    .C(_01234_),
    .D(_01239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01244_));
 sky130_fd_sc_hd__clkbuf_2 _06599_ (.A(_01196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01245_));
 sky130_fd_sc_hd__o21ai_1 _06600_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[23] ),
    .A2(_01242_),
    .B1(_01245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01246_));
 sky130_fd_sc_hd__nor2_1 _06601_ (.A(_01244_),
    .B(_01246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[23] ));
 sky130_fd_sc_hd__and2_1 _06602_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[24] ),
    .B(_01244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01247_));
 sky130_fd_sc_hd__o21ai_1 _06603_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[24] ),
    .A2(_01244_),
    .B1(_01245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01248_));
 sky130_fd_sc_hd__nor2_1 _06604_ (.A(_01247_),
    .B(_01248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[24] ));
 sky130_fd_sc_hd__o21ai_1 _06605_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[25] ),
    .A2(_01247_),
    .B1(_01245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01249_));
 sky130_fd_sc_hd__a21oi_1 _06606_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[25] ),
    .A2(_01247_),
    .B1(_01249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[25] ));
 sky130_fd_sc_hd__and4_1 _06607_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[24] ),
    .B(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[25] ),
    .C(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[26] ),
    .D(_01244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01250_));
 sky130_fd_sc_hd__a31o_1 _06608_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[24] ),
    .A2(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[25] ),
    .A3(_01244_),
    .B1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01251_));
 sky130_fd_sc_hd__and3b_1 _06609_ (.A_N(_01250_),
    .B(_01207_),
    .C(_01251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01252_));
 sky130_fd_sc_hd__clkbuf_1 _06610_ (.A(_01252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[26] ));
 sky130_fd_sc_hd__and2_1 _06611_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[27] ),
    .B(_01250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01253_));
 sky130_fd_sc_hd__o21ai_1 _06612_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[27] ),
    .A2(_01250_),
    .B1(_01245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01254_));
 sky130_fd_sc_hd__nor2_1 _06613_ (.A(_01253_),
    .B(_01254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[27] ));
 sky130_fd_sc_hd__and3_1 _06614_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[27] ),
    .B(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[28] ),
    .C(_01250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01255_));
 sky130_fd_sc_hd__o21ai_1 _06615_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[28] ),
    .A2(_01253_),
    .B1(_01245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01256_));
 sky130_fd_sc_hd__nor2_1 _06616_ (.A(_01255_),
    .B(_01256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[28] ));
 sky130_fd_sc_hd__o21ai_1 _06617_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[29] ),
    .A2(_01255_),
    .B1(_01207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01257_));
 sky130_fd_sc_hd__a21oi_1 _06618_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[29] ),
    .A2(_01255_),
    .B1(_01257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[29] ));
 sky130_fd_sc_hd__and3_1 _06619_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[28] ),
    .B(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[29] ),
    .C(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01258_));
 sky130_fd_sc_hd__and3_1 _06620_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[27] ),
    .B(_01250_),
    .C(_01258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01259_));
 sky130_fd_sc_hd__a21o_1 _06621_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[29] ),
    .A2(_01255_),
    .B1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01260_));
 sky130_fd_sc_hd__and3b_1 _06622_ (.A_N(_01259_),
    .B(_01058_),
    .C(_01260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01261_));
 sky130_fd_sc_hd__clkbuf_1 _06623_ (.A(_01261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[30] ));
 sky130_fd_sc_hd__o21ai_1 _06624_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[31] ),
    .A2(_01259_),
    .B1(_01207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01262_));
 sky130_fd_sc_hd__a21oi_1 _06625_ (.A1(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[31] ),
    .A2(_01259_),
    .B1(_01262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[31] ));
 sky130_fd_sc_hd__xor2_4 _06626_ (.A(\sa_inst._06_[10] ),
    .B(\sa_inst.sak._00_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01263_));
 sky130_fd_sc_hd__clkbuf_2 _06627_ (.A(_01263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01264_));
 sky130_fd_sc_hd__clkbuf_2 _06628_ (.A(_01264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._01_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06629_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._00_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01265_));
 sky130_fd_sc_hd__clkbuf_4 _06630_ (.A(_01265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01266_));
 sky130_fd_sc_hd__inv_2 _06631_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01267_));
 sky130_fd_sc_hd__clkbuf_2 _06632_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _06633_ (.A0(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ),
    .A1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[1] ),
    .S(_01268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01269_));
 sky130_fd_sc_hd__and2b_1 _06634_ (.A_N(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._22_ ),
    .B(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01270_));
 sky130_fd_sc_hd__mux4_2 _06635_ (.A0(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .A1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .A2(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .A3(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .S0(_01268_),
    .S1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01271_));
 sky130_fd_sc_hd__nor2_2 _06636_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._22_ ),
    .B(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01272_));
 sky130_fd_sc_hd__a32o_4 _06637_ (.A1(_01267_),
    .A2(_01269_),
    .A3(_01270_),
    .B1(_01271_),
    .B2(_01272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01273_));
 sky130_fd_sc_hd__xor2_4 _06638_ (.A(_01266_),
    .B(_01273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01274_));
 sky130_fd_sc_hd__buf_2 _06639_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01275_));
 sky130_fd_sc_hd__nand2_1 _06640_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[0] ),
    .B(_01275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01276_));
 sky130_fd_sc_hd__xnor2_1 _06641_ (.A(_01274_),
    .B(_01276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[0] ));
 sky130_fd_sc_hd__inv_2 _06642_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._22_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01277_));
 sky130_fd_sc_hd__clkbuf_2 _06643_ (.A(_01277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _06644_ (.A0(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .A1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .S(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _06645_ (.A0(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .A1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .S(_01268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _06646_ (.A0(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ),
    .A1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[2] ),
    .S(_01268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01281_));
 sky130_fd_sc_hd__clkbuf_2 _06647_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01282_));
 sky130_fd_sc_hd__and2b_1 _06648_ (.A_N(_01282_),
    .B(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01283_));
 sky130_fd_sc_hd__buf_2 _06649_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01284_));
 sky130_fd_sc_hd__clkbuf_2 _06650_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01285_));
 sky130_fd_sc_hd__mux4_2 _06651_ (.A0(_01279_),
    .A1(_01280_),
    .A2(_01281_),
    .A3(_01283_),
    .S0(_01284_),
    .S1(_01285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01286_));
 sky130_fd_sc_hd__nand4_4 _06652_ (.A(_01278_),
    .B(_01266_),
    .C(_01273_),
    .D(_01286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01287_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06653_ (.A(_01287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01288_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06654_ (.A(_01278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01289_));
 sky130_fd_sc_hd__a22o_1 _06655_ (.A1(_01266_),
    .A2(_01273_),
    .B1(_01286_),
    .B2(_01289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01290_));
 sky130_fd_sc_hd__and2_1 _06656_ (.A(_01288_),
    .B(_01290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01291_));
 sky130_fd_sc_hd__and3_1 _06657_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[1] ),
    .B(_01287_),
    .C(_01290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01292_));
 sky130_fd_sc_hd__a21oi_1 _06658_ (.A1(_01288_),
    .A2(_01290_),
    .B1(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01293_));
 sky130_fd_sc_hd__or2_1 _06659_ (.A(_01292_),
    .B(_01293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01294_));
 sky130_fd_sc_hd__nand2_1 _06660_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[0] ),
    .B(_01274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01295_));
 sky130_fd_sc_hd__xor2_1 _06661_ (.A(_01294_),
    .B(_01295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01296_));
 sky130_fd_sc_hd__buf_4 _06662_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _06663_ (.A0(_01291_),
    .A1(_01296_),
    .S(_01297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01298_));
 sky130_fd_sc_hd__clkbuf_1 _06664_ (.A(_01298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[1] ));
 sky130_fd_sc_hd__buf_2 _06665_ (.A(_01275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01299_));
 sky130_fd_sc_hd__o21ba_1 _06666_ (.A1(_01293_),
    .A2(_01295_),
    .B1_N(_01292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _06667_ (.A0(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._00_ ),
    .A1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .S(_01282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _06668_ (.A0(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .A1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .S(_01282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01302_));
 sky130_fd_sc_hd__clkbuf_2 _06669_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _06670_ (.A0(_01301_),
    .A1(_01302_),
    .S(_01303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01304_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06671_ (.A(_01267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _06672_ (.A0(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .A1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ),
    .S(_01282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01306_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06673_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01307_));
 sky130_fd_sc_hd__and3b_1 _06674_ (.A_N(_01307_),
    .B(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[1] ),
    .C(_01284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01308_));
 sky130_fd_sc_hd__a21o_1 _06675_ (.A1(_01305_),
    .A2(_01306_),
    .B1(_01308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01309_));
 sky130_fd_sc_hd__a22oi_4 _06676_ (.A1(_01272_),
    .A2(_01304_),
    .B1(_01309_),
    .B2(_01270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01310_));
 sky130_fd_sc_hd__xor2_1 _06677_ (.A(_01287_),
    .B(_01310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01311_));
 sky130_fd_sc_hd__nor2_1 _06678_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[2] ),
    .B(_01311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01312_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06679_ (.A(_01311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01313_));
 sky130_fd_sc_hd__and2_1 _06680_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[2] ),
    .B(_01313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01314_));
 sky130_fd_sc_hd__or3_1 _06681_ (.A(_01300_),
    .B(_01312_),
    .C(_01314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01315_));
 sky130_fd_sc_hd__o21ai_1 _06682_ (.A1(_01312_),
    .A2(_01314_),
    .B1(_01300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01316_));
 sky130_fd_sc_hd__clkinv_2 _06683_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01317_));
 sky130_fd_sc_hd__clkbuf_4 _06684_ (.A(_01317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01318_));
 sky130_fd_sc_hd__and2_1 _06685_ (.A(_01318_),
    .B(_01313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01319_));
 sky130_fd_sc_hd__a31o_1 _06686_ (.A1(_01299_),
    .A2(_01315_),
    .A3(_01316_),
    .B1(_01319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[2] ));
 sky130_fd_sc_hd__mux4_2 _06687_ (.A0(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._00_ ),
    .A1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .A2(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .A3(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .S0(_01284_),
    .S1(_01307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01320_));
 sky130_fd_sc_hd__mux4_1 _06688_ (.A0(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .A1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[2] ),
    .A2(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ),
    .A3(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[0] ),
    .S0(_01284_),
    .S1(_01307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01321_));
 sky130_fd_sc_hd__a22o_1 _06689_ (.A1(_01272_),
    .A2(_01320_),
    .B1(_01321_),
    .B2(_01270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01322_));
 sky130_fd_sc_hd__nor3b_2 _06690_ (.A(_01287_),
    .B(_01310_),
    .C_N(_01322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01323_));
 sky130_fd_sc_hd__clkbuf_2 _06691_ (.A(_01323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01324_));
 sky130_fd_sc_hd__o21bai_1 _06692_ (.A1(_01288_),
    .A2(_01310_),
    .B1_N(_01322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01325_));
 sky130_fd_sc_hd__and2b_1 _06693_ (.A_N(_01324_),
    .B(_01325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01326_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06694_ (.A(_01326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01327_));
 sky130_fd_sc_hd__nor2_1 _06695_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[3] ),
    .B(_01326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01328_));
 sky130_fd_sc_hd__nand3b_1 _06696_ (.A_N(_01324_),
    .B(_01325_),
    .C(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01329_));
 sky130_fd_sc_hd__or2b_1 _06697_ (.A(_01328_),
    .B_N(_01329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01330_));
 sky130_fd_sc_hd__nand2_1 _06698_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[2] ),
    .B(_01313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01331_));
 sky130_fd_sc_hd__o21ai_1 _06699_ (.A1(_01300_),
    .A2(_01312_),
    .B1(_01331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01332_));
 sky130_fd_sc_hd__xnor2_1 _06700_ (.A(_01330_),
    .B(_01332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01333_));
 sky130_fd_sc_hd__mux2_1 _06701_ (.A0(_01327_),
    .A1(_01333_),
    .S(_01297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01334_));
 sky130_fd_sc_hd__clkbuf_1 _06702_ (.A(_01334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[3] ));
 sky130_fd_sc_hd__clkbuf_2 _06703_ (.A(_01318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _06704_ (.A0(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .A1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .S(_01268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _06705_ (.A0(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .A1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .S(_01282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01337_));
 sky130_fd_sc_hd__mux4_1 _06706_ (.A0(_01265_),
    .A1(_01336_),
    .A2(_01337_),
    .A3(_01269_),
    .S0(_01284_),
    .S1(_01285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01338_));
 sky130_fd_sc_hd__nand2_1 _06707_ (.A(_01289_),
    .B(_01338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01339_));
 sky130_fd_sc_hd__xnor2_2 _06708_ (.A(_01323_),
    .B(_01339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01340_));
 sky130_fd_sc_hd__clkbuf_2 _06709_ (.A(_01340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01341_));
 sky130_fd_sc_hd__xnor2_1 _06710_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[4] ),
    .B(_01340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01342_));
 sky130_fd_sc_hd__o211a_1 _06711_ (.A1(_01300_),
    .A2(_01312_),
    .B1(_01331_),
    .C1(_01329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01343_));
 sky130_fd_sc_hd__or3_1 _06712_ (.A(_01328_),
    .B(_01342_),
    .C(_01343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01344_));
 sky130_fd_sc_hd__o21ai_1 _06713_ (.A1(_01328_),
    .A2(_01343_),
    .B1(_01342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01345_));
 sky130_fd_sc_hd__and3_1 _06714_ (.A(_01275_),
    .B(_01344_),
    .C(_01345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01346_));
 sky130_fd_sc_hd__a21o_1 _06715_ (.A1(_01335_),
    .A2(_01341_),
    .B1(_01346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[4] ));
 sky130_fd_sc_hd__inv_2 _06716_ (.A(_01339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01347_));
 sky130_fd_sc_hd__mux4_1 _06717_ (.A0(_01265_),
    .A1(_01279_),
    .A2(_01280_),
    .A3(_01281_),
    .S0(_01303_),
    .S1(_01285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01348_));
 sky130_fd_sc_hd__a22o_1 _06718_ (.A1(_01324_),
    .A2(_01347_),
    .B1(_01348_),
    .B2(_01289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01349_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06719_ (.A(_01324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01350_));
 sky130_fd_sc_hd__and3_1 _06720_ (.A(_01278_),
    .B(_01338_),
    .C(_01348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01351_));
 sky130_fd_sc_hd__nand2_2 _06721_ (.A(_01350_),
    .B(_01351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01352_));
 sky130_fd_sc_hd__and2_1 _06722_ (.A(_01349_),
    .B(_01352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01353_));
 sky130_fd_sc_hd__clkbuf_2 _06723_ (.A(_01353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01354_));
 sky130_fd_sc_hd__nand2_1 _06724_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[5] ),
    .B(_01354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01355_));
 sky130_fd_sc_hd__clkinv_2 _06725_ (.A(_01355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01356_));
 sky130_fd_sc_hd__nor2_1 _06726_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[5] ),
    .B(_01354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01357_));
 sky130_fd_sc_hd__or2_1 _06727_ (.A(_01356_),
    .B(_01357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01358_));
 sky130_fd_sc_hd__and2_1 _06728_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[4] ),
    .B(_01341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01359_));
 sky130_fd_sc_hd__inv_2 _06729_ (.A(_01359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01360_));
 sky130_fd_sc_hd__and2_1 _06730_ (.A(_01360_),
    .B(_01344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01361_));
 sky130_fd_sc_hd__xnor2_1 _06731_ (.A(_01358_),
    .B(_01361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01362_));
 sky130_fd_sc_hd__clkbuf_2 _06732_ (.A(_01317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01363_));
 sky130_fd_sc_hd__and3_1 _06733_ (.A(_01363_),
    .B(_01349_),
    .C(_01352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01364_));
 sky130_fd_sc_hd__o21bai_1 _06734_ (.A1(_01335_),
    .A2(_01362_),
    .B1_N(_01364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[5] ));
 sky130_fd_sc_hd__mux4_1 _06735_ (.A0(_01265_),
    .A1(_01301_),
    .A2(_01302_),
    .A3(_01306_),
    .S0(_01303_),
    .S1(_01285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01365_));
 sky130_fd_sc_hd__and2_2 _06736_ (.A(_01278_),
    .B(_01365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01366_));
 sky130_fd_sc_hd__xnor2_4 _06737_ (.A(_01352_),
    .B(_01366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01367_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06738_ (.A(_01367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01368_));
 sky130_fd_sc_hd__xnor2_1 _06739_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[6] ),
    .B(_01367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01369_));
 sky130_fd_sc_hd__a311o_1 _06740_ (.A1(_01360_),
    .A2(_01344_),
    .A3(_01355_),
    .B1(_01357_),
    .C1(_01369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01370_));
 sky130_fd_sc_hd__clkbuf_4 _06741_ (.A(_01317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01371_));
 sky130_fd_sc_hd__o211a_1 _06742_ (.A1(_01357_),
    .A2(_01361_),
    .B1(_01369_),
    .C1(_01355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01372_));
 sky130_fd_sc_hd__nor2_1 _06743_ (.A(_01371_),
    .B(_01372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01373_));
 sky130_fd_sc_hd__a22o_1 _06744_ (.A1(_01335_),
    .A2(_01368_),
    .B1(_01370_),
    .B2(_01373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[6] ));
 sky130_fd_sc_hd__clkbuf_2 _06745_ (.A(_01285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _06746_ (.A0(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._00_ ),
    .A1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .S(_01307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01375_));
 sky130_fd_sc_hd__nor2_1 _06747_ (.A(_01303_),
    .B(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._00_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01376_));
 sky130_fd_sc_hd__o21ba_1 _06748_ (.A1(_01305_),
    .A2(_01375_),
    .B1_N(_01376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01377_));
 sky130_fd_sc_hd__inv_2 _06749_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01378_));
 sky130_fd_sc_hd__mux4_1 _06750_ (.A0(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .A1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .A2(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .A3(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ),
    .S0(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .S1(_01307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01379_));
 sky130_fd_sc_hd__or2_1 _06751_ (.A(_01378_),
    .B(_01379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01380_));
 sky130_fd_sc_hd__o211a_1 _06752_ (.A1(_01374_),
    .A2(_01377_),
    .B1(_01380_),
    .C1(_01278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01381_));
 sky130_fd_sc_hd__and3_1 _06753_ (.A(_01351_),
    .B(_01366_),
    .C(_01381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01382_));
 sky130_fd_sc_hd__nand2_1 _06754_ (.A(_01350_),
    .B(_01382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01383_));
 sky130_fd_sc_hd__a31o_1 _06755_ (.A1(_01350_),
    .A2(_01351_),
    .A3(_01366_),
    .B1(_01381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01384_));
 sky130_fd_sc_hd__and2_1 _06756_ (.A(_01383_),
    .B(_01384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01385_));
 sky130_fd_sc_hd__nor2_1 _06757_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[7] ),
    .B(_01385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01386_));
 sky130_fd_sc_hd__and3_1 _06758_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[7] ),
    .B(_01383_),
    .C(_01384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01387_));
 sky130_fd_sc_hd__or2_1 _06759_ (.A(_01386_),
    .B(_01387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01388_));
 sky130_fd_sc_hd__and2_1 _06760_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[6] ),
    .B(_01368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01389_));
 sky130_fd_sc_hd__or2b_1 _06761_ (.A(_01389_),
    .B_N(_01370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01390_));
 sky130_fd_sc_hd__xnor2_1 _06762_ (.A(_01388_),
    .B(_01390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01391_));
 sky130_fd_sc_hd__clkbuf_2 _06763_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01392_));
 sky130_fd_sc_hd__buf_2 _06764_ (.A(_01392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _06765_ (.A0(_01385_),
    .A1(_01391_),
    .S(_01393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01394_));
 sky130_fd_sc_hd__clkbuf_1 _06766_ (.A(_01394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[7] ));
 sky130_fd_sc_hd__or2_1 _06767_ (.A(_01378_),
    .B(_01271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01395_));
 sky130_fd_sc_hd__o21a_1 _06768_ (.A1(_01374_),
    .A2(_01265_),
    .B1(_01277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01396_));
 sky130_fd_sc_hd__and2_1 _06769_ (.A(_01395_),
    .B(_01396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01397_));
 sky130_fd_sc_hd__nand3_1 _06770_ (.A(_01350_),
    .B(_01382_),
    .C(_01397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01398_));
 sky130_fd_sc_hd__a21o_1 _06771_ (.A1(_01324_),
    .A2(_01382_),
    .B1(_01397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01399_));
 sky130_fd_sc_hd__and2_1 _06772_ (.A(_01398_),
    .B(_01399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01400_));
 sky130_fd_sc_hd__clkbuf_2 _06773_ (.A(_01400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01401_));
 sky130_fd_sc_hd__xnor2_1 _06774_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[8] ),
    .B(_01401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01402_));
 sky130_fd_sc_hd__nor2_1 _06775_ (.A(_01389_),
    .B(_01387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01403_));
 sky130_fd_sc_hd__a21o_1 _06776_ (.A1(_01370_),
    .A2(_01403_),
    .B1(_01386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01404_));
 sky130_fd_sc_hd__or2_1 _06777_ (.A(_01402_),
    .B(_01404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01405_));
 sky130_fd_sc_hd__a21oi_1 _06778_ (.A1(_01402_),
    .A2(_01404_),
    .B1(_01371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01406_));
 sky130_fd_sc_hd__a22o_1 _06779_ (.A1(_01335_),
    .A2(_01401_),
    .B1(_01405_),
    .B2(_01406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[8] ));
 sky130_fd_sc_hd__clkbuf_4 _06780_ (.A(_01392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01407_));
 sky130_fd_sc_hd__nand2_1 _06781_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[8] ),
    .B(_01401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01408_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06782_ (.A(_01378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _06783_ (.A0(_01279_),
    .A1(_01280_),
    .S(_01303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01410_));
 sky130_fd_sc_hd__o21a_1 _06784_ (.A1(_01409_),
    .A2(_01410_),
    .B1(_01396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01411_));
 sky130_fd_sc_hd__and2_1 _06785_ (.A(_01395_),
    .B(_01411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01412_));
 sky130_fd_sc_hd__nand3_1 _06786_ (.A(_01323_),
    .B(_01382_),
    .C(_01412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01413_));
 sky130_fd_sc_hd__buf_2 _06787_ (.A(_01413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01414_));
 sky130_fd_sc_hd__a31o_2 _06788_ (.A1(_01350_),
    .A2(_01382_),
    .A3(_01397_),
    .B1(_01411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01415_));
 sky130_fd_sc_hd__and3_1 _06789_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[9] ),
    .B(_01414_),
    .C(_01415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01416_));
 sky130_fd_sc_hd__a21oi_1 _06790_ (.A1(_01414_),
    .A2(_01415_),
    .B1(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01417_));
 sky130_fd_sc_hd__or2_1 _06791_ (.A(_01416_),
    .B(_01417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01418_));
 sky130_fd_sc_hd__a21o_1 _06792_ (.A1(_01408_),
    .A2(_01405_),
    .B1(_01418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01419_));
 sky130_fd_sc_hd__nand2_1 _06793_ (.A(_01407_),
    .B(_01419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01420_));
 sky130_fd_sc_hd__and3_1 _06794_ (.A(_01408_),
    .B(_01405_),
    .C(_01418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01421_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06795_ (.A(_01414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01422_));
 sky130_fd_sc_hd__and2_1 _06796_ (.A(_01422_),
    .B(_01415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01423_));
 sky130_fd_sc_hd__a2bb2o_1 _06797_ (.A1_N(_01420_),
    .A2_N(_01421_),
    .B1(_01423_),
    .B2(_01335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[9] ));
 sky130_fd_sc_hd__o21ai_2 _06798_ (.A1(_01374_),
    .A2(_01266_),
    .B1(_01289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01424_));
 sky130_fd_sc_hd__nor2_1 _06799_ (.A(_01409_),
    .B(_01304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01425_));
 sky130_fd_sc_hd__nor2_1 _06800_ (.A(_01424_),
    .B(_01425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01426_));
 sky130_fd_sc_hd__xnor2_1 _06801_ (.A(_01413_),
    .B(_01426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01427_));
 sky130_fd_sc_hd__xnor2_1 _06802_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[10] ),
    .B(_01427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01428_));
 sky130_fd_sc_hd__a21oi_1 _06803_ (.A1(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[8] ),
    .A2(_01401_),
    .B1(_01416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01429_));
 sky130_fd_sc_hd__a21o_1 _06804_ (.A1(_01405_),
    .A2(_01429_),
    .B1(_01417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01430_));
 sky130_fd_sc_hd__or2_1 _06805_ (.A(_01428_),
    .B(_01430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01431_));
 sky130_fd_sc_hd__nand2_1 _06806_ (.A(_01428_),
    .B(_01430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01432_));
 sky130_fd_sc_hd__clkbuf_2 _06807_ (.A(_01427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01433_));
 sky130_fd_sc_hd__and2_1 _06808_ (.A(_01363_),
    .B(_01433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01434_));
 sky130_fd_sc_hd__a31o_1 _06809_ (.A1(_01299_),
    .A2(_01431_),
    .A3(_01432_),
    .B1(_01434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[10] ));
 sky130_fd_sc_hd__nand2_1 _06810_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[10] ),
    .B(_01433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01435_));
 sky130_fd_sc_hd__inv_2 _06811_ (.A(_01426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01436_));
 sky130_fd_sc_hd__nor2_2 _06812_ (.A(_01409_),
    .B(_01320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01437_));
 sky130_fd_sc_hd__or3_1 _06813_ (.A(_01413_),
    .B(_01436_),
    .C(_01437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01438_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06814_ (.A(_01438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01439_));
 sky130_fd_sc_hd__o22ai_4 _06815_ (.A1(_01414_),
    .A2(_01436_),
    .B1(_01437_),
    .B2(_01424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01440_));
 sky130_fd_sc_hd__and3_1 _06816_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[11] ),
    .B(_01439_),
    .C(_01440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01441_));
 sky130_fd_sc_hd__a21oi_1 _06817_ (.A1(_01439_),
    .A2(_01440_),
    .B1(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01442_));
 sky130_fd_sc_hd__or2_1 _06818_ (.A(_01441_),
    .B(_01442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01443_));
 sky130_fd_sc_hd__a21o_1 _06819_ (.A1(_01435_),
    .A2(_01431_),
    .B1(_01443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01444_));
 sky130_fd_sc_hd__nand3_1 _06820_ (.A(_01435_),
    .B(_01431_),
    .C(_01443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01445_));
 sky130_fd_sc_hd__and3_1 _06821_ (.A(_01363_),
    .B(_01439_),
    .C(_01440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01446_));
 sky130_fd_sc_hd__a31o_1 _06822_ (.A1(_01299_),
    .A2(_01444_),
    .A3(_01445_),
    .B1(_01446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[11] ));
 sky130_fd_sc_hd__a21o_1 _06823_ (.A1(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[10] ),
    .A2(_01433_),
    .B1(_01441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01447_));
 sky130_fd_sc_hd__or2b_1 _06824_ (.A(_01442_),
    .B_N(_01447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01448_));
 sky130_fd_sc_hd__or3_1 _06825_ (.A(_01428_),
    .B(_01441_),
    .C(_01442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01449_));
 sky130_fd_sc_hd__or3_1 _06826_ (.A(_01417_),
    .B(_01429_),
    .C(_01449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01450_));
 sky130_fd_sc_hd__or2_1 _06827_ (.A(_01402_),
    .B(_01418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01451_));
 sky130_fd_sc_hd__a2111o_1 _06828_ (.A1(_01370_),
    .A2(_01403_),
    .B1(_01449_),
    .C1(_01451_),
    .D1(_01386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01452_));
 sky130_fd_sc_hd__o21ba_1 _06829_ (.A1(_01305_),
    .A2(_01336_),
    .B1_N(_01376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01453_));
 sky130_fd_sc_hd__o31a_2 _06830_ (.A1(_01422_),
    .A2(_01425_),
    .A3(_01437_),
    .B1(_01396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01454_));
 sky130_fd_sc_hd__o21a_2 _06831_ (.A1(_01409_),
    .A2(_01453_),
    .B1(_01454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01455_));
 sky130_fd_sc_hd__nand2_1 _06832_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[12] ),
    .B(_01455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01456_));
 sky130_fd_sc_hd__or2_1 _06833_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[12] ),
    .B(_01455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01457_));
 sky130_fd_sc_hd__nand2_1 _06834_ (.A(_01456_),
    .B(_01457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01458_));
 sky130_fd_sc_hd__a31o_1 _06835_ (.A1(_01448_),
    .A2(_01450_),
    .A3(_01452_),
    .B1(_01458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01459_));
 sky130_fd_sc_hd__clkbuf_4 _06836_ (.A(_01317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01460_));
 sky130_fd_sc_hd__a41oi_1 _06837_ (.A1(_01458_),
    .A2(_01448_),
    .A3(_01450_),
    .A4(_01452_),
    .B1(_01460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01461_));
 sky130_fd_sc_hd__and2_1 _06838_ (.A(_01318_),
    .B(_01455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01462_));
 sky130_fd_sc_hd__a21o_1 _06839_ (.A1(_01459_),
    .A2(_01461_),
    .B1(_01462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[12] ));
 sky130_fd_sc_hd__clkbuf_1 _06840_ (.A(_01454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01463_));
 sky130_fd_sc_hd__nor2_1 _06841_ (.A(_01305_),
    .B(_01279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01464_));
 sky130_fd_sc_hd__o21ai_2 _06842_ (.A1(_01376_),
    .A2(_01464_),
    .B1(_01374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01465_));
 sky130_fd_sc_hd__clkbuf_1 _06843_ (.A(_01465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01466_));
 sky130_fd_sc_hd__and3_1 _06844_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[13] ),
    .B(_01463_),
    .C(_01466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01467_));
 sky130_fd_sc_hd__a21oi_1 _06845_ (.A1(_01454_),
    .A2(_01465_),
    .B1(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01468_));
 sky130_fd_sc_hd__nand2_1 _06846_ (.A(_01456_),
    .B(_01459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01469_));
 sky130_fd_sc_hd__o21bai_1 _06847_ (.A1(_01467_),
    .A2(_01468_),
    .B1_N(_01469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01470_));
 sky130_fd_sc_hd__or3b_1 _06848_ (.A(_01467_),
    .B(_01468_),
    .C_N(_01469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01471_));
 sky130_fd_sc_hd__and3_1 _06849_ (.A(_01363_),
    .B(_01463_),
    .C(_01466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01472_));
 sky130_fd_sc_hd__a31o_1 _06850_ (.A1(_01299_),
    .A2(_01470_),
    .A3(_01471_),
    .B1(_01472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[13] ));
 sky130_fd_sc_hd__nor2_1 _06851_ (.A(_01467_),
    .B(_01469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01473_));
 sky130_fd_sc_hd__nor2_1 _06852_ (.A(_01305_),
    .B(_01301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01474_));
 sky130_fd_sc_hd__o21ai_1 _06853_ (.A1(_01376_),
    .A2(_01474_),
    .B1(_01374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01475_));
 sky130_fd_sc_hd__o311a_2 _06854_ (.A1(_01422_),
    .A2(_01425_),
    .A3(_01437_),
    .B1(_01475_),
    .C1(_01396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01476_));
 sky130_fd_sc_hd__xnor2_1 _06855_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[14] ),
    .B(_01476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01477_));
 sky130_fd_sc_hd__o21ai_1 _06856_ (.A1(_01468_),
    .A2(_01473_),
    .B1(_01477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01478_));
 sky130_fd_sc_hd__or2_1 _06857_ (.A(_01468_),
    .B(_01477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01479_));
 sky130_fd_sc_hd__or2_1 _06858_ (.A(_01473_),
    .B(_01479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01480_));
 sky130_fd_sc_hd__and2_1 _06859_ (.A(_01318_),
    .B(_01476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01481_));
 sky130_fd_sc_hd__a31o_1 _06860_ (.A1(_01299_),
    .A2(_01478_),
    .A3(_01480_),
    .B1(_01481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[14] ));
 sky130_fd_sc_hd__clkbuf_2 _06861_ (.A(_01275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01482_));
 sky130_fd_sc_hd__nand2_1 _06862_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[14] ),
    .B(_01476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01483_));
 sky130_fd_sc_hd__or2_1 _06863_ (.A(_01409_),
    .B(_01377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01484_));
 sky130_fd_sc_hd__o311a_1 _06864_ (.A1(_01422_),
    .A2(_01425_),
    .A3(_01437_),
    .B1(_01484_),
    .C1(_01396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01485_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06865_ (.A(_01485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01486_));
 sky130_fd_sc_hd__nand2_1 _06866_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[15] ),
    .B(_01486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01487_));
 sky130_fd_sc_hd__or2_1 _06867_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[15] ),
    .B(_01486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01488_));
 sky130_fd_sc_hd__nand2_1 _06868_ (.A(_01487_),
    .B(_01488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01489_));
 sky130_fd_sc_hd__a21o_1 _06869_ (.A1(_01483_),
    .A2(_01480_),
    .B1(_01489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01490_));
 sky130_fd_sc_hd__nand3_1 _06870_ (.A(_01483_),
    .B(_01480_),
    .C(_01489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01491_));
 sky130_fd_sc_hd__and2_1 _06871_ (.A(_01363_),
    .B(_01486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01492_));
 sky130_fd_sc_hd__a31o_1 _06872_ (.A1(_01482_),
    .A2(_01490_),
    .A3(_01491_),
    .B1(_01492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[15] ));
 sky130_fd_sc_hd__buf_2 _06873_ (.A(_01392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01493_));
 sky130_fd_sc_hd__clkbuf_4 _06874_ (.A(_01493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01494_));
 sky130_fd_sc_hd__nand3_1 _06875_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[13] ),
    .B(_01463_),
    .C(_01466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01495_));
 sky130_fd_sc_hd__nor2_1 _06876_ (.A(_01479_),
    .B(_01489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01496_));
 sky130_fd_sc_hd__nand2_1 _06877_ (.A(_01495_),
    .B(_01496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01497_));
 sky130_fd_sc_hd__a21bo_1 _06878_ (.A1(_01483_),
    .A2(_01487_),
    .B1_N(_01488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01498_));
 sky130_fd_sc_hd__a211o_1 _06879_ (.A1(_01456_),
    .A2(_01495_),
    .B1(_01479_),
    .C1(_01489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01499_));
 sky130_fd_sc_hd__o211ai_4 _06880_ (.A1(_01459_),
    .A2(_01497_),
    .B1(_01498_),
    .C1(_01499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01500_));
 sky130_fd_sc_hd__and3_1 _06881_ (.A(_01289_),
    .B(_01266_),
    .C(_01438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01501_));
 sky130_fd_sc_hd__clkbuf_2 _06882_ (.A(_01501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01502_));
 sky130_fd_sc_hd__clkbuf_2 _06883_ (.A(_01502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01503_));
 sky130_fd_sc_hd__nand2_1 _06884_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[16] ),
    .B(_01503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01504_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06885_ (.A(_01501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01505_));
 sky130_fd_sc_hd__or2_1 _06886_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[16] ),
    .B(_01505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01506_));
 sky130_fd_sc_hd__nand2_1 _06887_ (.A(_01504_),
    .B(_01506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01507_));
 sky130_fd_sc_hd__xnor2_1 _06888_ (.A(_01500_),
    .B(_01507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01508_));
 sky130_fd_sc_hd__buf_2 _06889_ (.A(_01502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01509_));
 sky130_fd_sc_hd__clkbuf_2 _06890_ (.A(_01509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01510_));
 sky130_fd_sc_hd__clkbuf_2 _06891_ (.A(_01510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01511_));
 sky130_fd_sc_hd__clkbuf_2 _06892_ (.A(_01511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01512_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06893_ (.A(_01512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01513_));
 sky130_fd_sc_hd__clkbuf_2 _06894_ (.A(_01513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01514_));
 sky130_fd_sc_hd__and2_1 _06895_ (.A(_01317_),
    .B(_01514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01515_));
 sky130_fd_sc_hd__buf_2 _06896_ (.A(_01515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01516_));
 sky130_fd_sc_hd__clkbuf_2 _06897_ (.A(_01516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01517_));
 sky130_fd_sc_hd__a21o_1 _06898_ (.A1(_01494_),
    .A2(_01508_),
    .B1(_01517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[16] ));
 sky130_fd_sc_hd__inv_2 _06899_ (.A(_01500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01518_));
 sky130_fd_sc_hd__o21a_1 _06900_ (.A1(_01518_),
    .A2(_01507_),
    .B1(_01504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01519_));
 sky130_fd_sc_hd__nand2_1 _06901_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[17] ),
    .B(_01509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01520_));
 sky130_fd_sc_hd__clkbuf_2 _06902_ (.A(_01502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01521_));
 sky130_fd_sc_hd__or2_1 _06903_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[17] ),
    .B(_01521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01522_));
 sky130_fd_sc_hd__nand2_1 _06904_ (.A(_01520_),
    .B(_01522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01523_));
 sky130_fd_sc_hd__or2_1 _06905_ (.A(_01519_),
    .B(_01523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01524_));
 sky130_fd_sc_hd__nand2_1 _06906_ (.A(_01519_),
    .B(_01523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01525_));
 sky130_fd_sc_hd__clkbuf_2 _06907_ (.A(_01516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01526_));
 sky130_fd_sc_hd__a31o_1 _06908_ (.A1(_01482_),
    .A2(_01524_),
    .A3(_01525_),
    .B1(_01526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[17] ));
 sky130_fd_sc_hd__or2b_1 _06909_ (.A(_01519_),
    .B_N(_01522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01527_));
 sky130_fd_sc_hd__nand2_1 _06910_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[18] ),
    .B(_01509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01528_));
 sky130_fd_sc_hd__or2_1 _06911_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[18] ),
    .B(_01521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01529_));
 sky130_fd_sc_hd__nand2_1 _06912_ (.A(_01528_),
    .B(_01529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01530_));
 sky130_fd_sc_hd__a21o_1 _06913_ (.A1(_01520_),
    .A2(_01527_),
    .B1(_01530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01531_));
 sky130_fd_sc_hd__nand3_1 _06914_ (.A(_01520_),
    .B(_01527_),
    .C(_01530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01532_));
 sky130_fd_sc_hd__a31o_1 _06915_ (.A1(_01482_),
    .A2(_01531_),
    .A3(_01532_),
    .B1(_01526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[18] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06916_ (.A(_01505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01533_));
 sky130_fd_sc_hd__xnor2_1 _06917_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[19] ),
    .B(_01533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01534_));
 sky130_fd_sc_hd__a21o_1 _06918_ (.A1(_01528_),
    .A2(_01531_),
    .B1(_01534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01535_));
 sky130_fd_sc_hd__nand3_1 _06919_ (.A(_01528_),
    .B(_01531_),
    .C(_01534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01536_));
 sky130_fd_sc_hd__a31o_1 _06920_ (.A1(_01482_),
    .A2(_01535_),
    .A3(_01536_),
    .B1(_01526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[19] ));
 sky130_fd_sc_hd__and2_1 _06921_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[20] ),
    .B(_01533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01537_));
 sky130_fd_sc_hd__nor2_1 _06922_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[20] ),
    .B(_01510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01538_));
 sky130_fd_sc_hd__or2_1 _06923_ (.A(_01537_),
    .B(_01538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01539_));
 sky130_fd_sc_hd__or4_1 _06924_ (.A(_01507_),
    .B(_01523_),
    .C(_01530_),
    .D(_01534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01540_));
 sky130_fd_sc_hd__buf_2 _06925_ (.A(_01511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01541_));
 sky130_fd_sc_hd__o41a_1 _06926_ (.A1(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[16] ),
    .A2(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[17] ),
    .A3(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[18] ),
    .A4(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[19] ),
    .B1(_01541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01542_));
 sky130_fd_sc_hd__o21ba_1 _06927_ (.A1(_01518_),
    .A2(_01540_),
    .B1_N(_01542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01543_));
 sky130_fd_sc_hd__nor2_1 _06928_ (.A(_01539_),
    .B(_01543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01544_));
 sky130_fd_sc_hd__a21o_1 _06929_ (.A1(_01539_),
    .A2(_01543_),
    .B1(_01460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01545_));
 sky130_fd_sc_hd__buf_2 _06930_ (.A(_01515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01546_));
 sky130_fd_sc_hd__o21bai_1 _06931_ (.A1(_01544_),
    .A2(_01545_),
    .B1_N(_01546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[20] ));
 sky130_fd_sc_hd__or2_1 _06932_ (.A(_01537_),
    .B(_01544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01547_));
 sky130_fd_sc_hd__and2_1 _06933_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[21] ),
    .B(_01533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01548_));
 sky130_fd_sc_hd__or2_1 _06934_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[21] ),
    .B(_01533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01549_));
 sky130_fd_sc_hd__or2b_1 _06935_ (.A(_01548_),
    .B_N(_01549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01550_));
 sky130_fd_sc_hd__xnor2_1 _06936_ (.A(_01547_),
    .B(_01550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01551_));
 sky130_fd_sc_hd__a21o_1 _06937_ (.A1(_01494_),
    .A2(_01551_),
    .B1(_01517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[21] ));
 sky130_fd_sc_hd__and2_1 _06938_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[22] ),
    .B(_01533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01552_));
 sky130_fd_sc_hd__nor2_1 _06939_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[22] ),
    .B(_01510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01553_));
 sky130_fd_sc_hd__nor2_1 _06940_ (.A(_01552_),
    .B(_01553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01554_));
 sky130_fd_sc_hd__o311a_1 _06941_ (.A1(_01537_),
    .A2(_01544_),
    .A3(_01548_),
    .B1(_01549_),
    .C1(_01554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01555_));
 sky130_fd_sc_hd__inv_2 _06942_ (.A(_01555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01556_));
 sky130_fd_sc_hd__a211o_1 _06943_ (.A1(_01547_),
    .A2(_01549_),
    .B1(_01554_),
    .C1(_01548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01557_));
 sky130_fd_sc_hd__a31o_1 _06944_ (.A1(_01482_),
    .A2(_01556_),
    .A3(_01557_),
    .B1(_01526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[22] ));
 sky130_fd_sc_hd__buf_2 _06945_ (.A(_01297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01558_));
 sky130_fd_sc_hd__xor2_1 _06946_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[23] ),
    .B(_01510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01559_));
 sky130_fd_sc_hd__o21ai_1 _06947_ (.A1(_01552_),
    .A2(_01555_),
    .B1(_01559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01560_));
 sky130_fd_sc_hd__or3_1 _06948_ (.A(_01552_),
    .B(_01555_),
    .C(_01559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01561_));
 sky130_fd_sc_hd__a31o_1 _06949_ (.A1(_01558_),
    .A2(_01560_),
    .A3(_01561_),
    .B1(_01526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[23] ));
 sky130_fd_sc_hd__nand2_1 _06950_ (.A(_01554_),
    .B(_01559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01562_));
 sky130_fd_sc_hd__nor4_1 _06951_ (.A(_01539_),
    .B(_01540_),
    .C(_01550_),
    .D(_01562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01563_));
 sky130_fd_sc_hd__o41a_1 _06952_ (.A1(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[20] ),
    .A2(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[21] ),
    .A3(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[22] ),
    .A4(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[23] ),
    .B1(_01541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01564_));
 sky130_fd_sc_hd__a211o_2 _06953_ (.A1(_01500_),
    .A2(_01563_),
    .B1(_01564_),
    .C1(_01542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01565_));
 sky130_fd_sc_hd__buf_2 _06954_ (.A(_01510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01566_));
 sky130_fd_sc_hd__xor2_1 _06955_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[24] ),
    .B(_01566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01567_));
 sky130_fd_sc_hd__nand2_1 _06956_ (.A(_01565_),
    .B(_01567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01568_));
 sky130_fd_sc_hd__o21a_1 _06957_ (.A1(_01565_),
    .A2(_01567_),
    .B1(_01493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01569_));
 sky130_fd_sc_hd__a21o_1 _06958_ (.A1(_01568_),
    .A2(_01569_),
    .B1(_01517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[24] ));
 sky130_fd_sc_hd__xor2_1 _06959_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[25] ),
    .B(_01566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01570_));
 sky130_fd_sc_hd__clkbuf_2 _06960_ (.A(_01541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01571_));
 sky130_fd_sc_hd__clkbuf_1 _06961_ (.A(_01571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01572_));
 sky130_fd_sc_hd__clkbuf_2 _06962_ (.A(_01572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01573_));
 sky130_fd_sc_hd__a22o_1 _06963_ (.A1(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[24] ),
    .A2(_01573_),
    .B1(_01565_),
    .B2(_01567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01574_));
 sky130_fd_sc_hd__xor2_1 _06964_ (.A(_01570_),
    .B(_01574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01575_));
 sky130_fd_sc_hd__a21o_1 _06965_ (.A1(_01494_),
    .A2(_01575_),
    .B1(_01517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[25] ));
 sky130_fd_sc_hd__o21ai_1 _06966_ (.A1(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[24] ),
    .A2(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[25] ),
    .B1(_01514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01576_));
 sky130_fd_sc_hd__and2_1 _06967_ (.A(_01567_),
    .B(_01570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01577_));
 sky130_fd_sc_hd__nand2_1 _06968_ (.A(_01565_),
    .B(_01577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01578_));
 sky130_fd_sc_hd__nand2_1 _06969_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[26] ),
    .B(_01541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01579_));
 sky130_fd_sc_hd__or2_1 _06970_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[26] ),
    .B(_01511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01580_));
 sky130_fd_sc_hd__nand2_1 _06971_ (.A(_01579_),
    .B(_01580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01581_));
 sky130_fd_sc_hd__a21o_1 _06972_ (.A1(_01576_),
    .A2(_01578_),
    .B1(_01581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01582_));
 sky130_fd_sc_hd__nand3_1 _06973_ (.A(_01581_),
    .B(_01576_),
    .C(_01578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01583_));
 sky130_fd_sc_hd__buf_2 _06974_ (.A(_01515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01584_));
 sky130_fd_sc_hd__a31o_1 _06975_ (.A1(_01558_),
    .A2(_01582_),
    .A3(_01583_),
    .B1(_01584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[26] ));
 sky130_fd_sc_hd__clkbuf_4 _06976_ (.A(_01493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01585_));
 sky130_fd_sc_hd__xnor2_1 _06977_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[27] ),
    .B(_01512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01586_));
 sky130_fd_sc_hd__nand2_1 _06978_ (.A(_01579_),
    .B(_01582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01587_));
 sky130_fd_sc_hd__xnor2_1 _06979_ (.A(_01586_),
    .B(_01587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01588_));
 sky130_fd_sc_hd__a21o_1 _06980_ (.A1(_01585_),
    .A2(_01588_),
    .B1(_01517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[27] ));
 sky130_fd_sc_hd__nor2_1 _06981_ (.A(_01581_),
    .B(_01586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01589_));
 sky130_fd_sc_hd__o41a_1 _06982_ (.A1(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[24] ),
    .A2(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[25] ),
    .A3(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[26] ),
    .A4(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[27] ),
    .B1(_01571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01590_));
 sky130_fd_sc_hd__a31oi_2 _06983_ (.A1(_01565_),
    .A2(_01577_),
    .A3(_01589_),
    .B1(_01590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01591_));
 sky130_fd_sc_hd__and2_1 _06984_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[28] ),
    .B(_01512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01592_));
 sky130_fd_sc_hd__nor2_1 _06985_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[28] ),
    .B(_01571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01593_));
 sky130_fd_sc_hd__or2_1 _06986_ (.A(_01592_),
    .B(_01593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01594_));
 sky130_fd_sc_hd__nor2_1 _06987_ (.A(_01591_),
    .B(_01594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01595_));
 sky130_fd_sc_hd__a21o_1 _06988_ (.A1(_01591_),
    .A2(_01594_),
    .B1(_01460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01596_));
 sky130_fd_sc_hd__o21bai_1 _06989_ (.A1(_01595_),
    .A2(_01596_),
    .B1_N(_01546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[28] ));
 sky130_fd_sc_hd__nand2_1 _06990_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[29] ),
    .B(_01513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01597_));
 sky130_fd_sc_hd__or2_1 _06991_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[29] ),
    .B(_01513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01598_));
 sky130_fd_sc_hd__o211ai_1 _06992_ (.A1(_01592_),
    .A2(_01595_),
    .B1(_01597_),
    .C1(_01598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01599_));
 sky130_fd_sc_hd__a211o_1 _06993_ (.A1(_01597_),
    .A2(_01598_),
    .B1(_01592_),
    .C1(_01595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01600_));
 sky130_fd_sc_hd__a31o_1 _06994_ (.A1(_01558_),
    .A2(_01599_),
    .A3(_01600_),
    .B1(_01584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[29] ));
 sky130_fd_sc_hd__o21ai_1 _06995_ (.A1(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[28] ),
    .A2(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[29] ),
    .B1(_01514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01601_));
 sky130_fd_sc_hd__or4bb_1 _06996_ (.A(_01591_),
    .B(_01594_),
    .C_N(_01597_),
    .D_N(_01598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01602_));
 sky130_fd_sc_hd__and2_1 _06997_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[30] ),
    .B(_01572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01603_));
 sky130_fd_sc_hd__nor2_1 _06998_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[30] ),
    .B(_01572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01604_));
 sky130_fd_sc_hd__or2_1 _06999_ (.A(_01603_),
    .B(_01604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01605_));
 sky130_fd_sc_hd__a21o_1 _07000_ (.A1(_01601_),
    .A2(_01602_),
    .B1(_01605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01606_));
 sky130_fd_sc_hd__nand3_1 _07001_ (.A(_01605_),
    .B(_01601_),
    .C(_01602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01607_));
 sky130_fd_sc_hd__a31o_1 _07002_ (.A1(_01558_),
    .A2(_01606_),
    .A3(_01607_),
    .B1(_01584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[30] ));
 sky130_fd_sc_hd__nand2_1 _07003_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[31] ),
    .B(_01573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01608_));
 sky130_fd_sc_hd__or2_1 _07004_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[31] ),
    .B(_01573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01609_));
 sky130_fd_sc_hd__a21oi_1 _07005_ (.A1(_01601_),
    .A2(_01602_),
    .B1(_01605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01610_));
 sky130_fd_sc_hd__a211o_1 _07006_ (.A1(_01608_),
    .A2(_01609_),
    .B1(_01603_),
    .C1(_01610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01611_));
 sky130_fd_sc_hd__o211ai_1 _07007_ (.A1(_01603_),
    .A2(_01610_),
    .B1(_01608_),
    .C1(_01609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01612_));
 sky130_fd_sc_hd__a31o_1 _07008_ (.A1(_01558_),
    .A2(_01611_),
    .A3(_01612_),
    .B1(_01584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[31] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07009_ (.A(\sa_inst.sak._00_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01613_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07010_ (.A(_01613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01614_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07011_ (.A(\sa_inst._06_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01615_));
 sky130_fd_sc_hd__nand2_1 _07012_ (.A(_01614_),
    .B(_01615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01616_));
 sky130_fd_sc_hd__xnor2_1 _07013_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._01_ ),
    .B(_01616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01617_));
 sky130_fd_sc_hd__clkbuf_2 _07014_ (.A(\sa_inst._06_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01618_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07015_ (.A(\sa_inst.sak._00_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01619_));
 sky130_fd_sc_hd__a22oi_1 _07016_ (.A1(_01614_),
    .A2(_01618_),
    .B1(_01619_),
    .B2(_01615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01620_));
 sky130_fd_sc_hd__and2_1 _07017_ (.A(\sa_inst._06_[5] ),
    .B(_01619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01621_));
 sky130_fd_sc_hd__and3_1 _07018_ (.A(_01614_),
    .B(_01615_),
    .C(_01621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01622_));
 sky130_fd_sc_hd__or2_1 _07019_ (.A(_01620_),
    .B(_01622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01623_));
 sky130_fd_sc_hd__xnor2_1 _07020_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._01_ ),
    .B(_01623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01624_));
 sky130_fd_sc_hd__xor2_4 _07021_ (.A(_01132_),
    .B(\sa_inst._06_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01625_));
 sky130_fd_sc_hd__clkbuf_2 _07022_ (.A(_01625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01626_));
 sky130_fd_sc_hd__mux2_1 _07023_ (.A0(_01617_),
    .A1(_01624_),
    .S(_01626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01627_));
 sky130_fd_sc_hd__clkbuf_1 _07024_ (.A(_01627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[1] ));
 sky130_fd_sc_hd__clkbuf_2 _07025_ (.A(\sa_inst._06_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01628_));
 sky130_fd_sc_hd__and3_1 _07026_ (.A(_01613_),
    .B(_01628_),
    .C(_01621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01629_));
 sky130_fd_sc_hd__a21oi_1 _07027_ (.A1(_01614_),
    .A2(_01628_),
    .B1(_01621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01630_));
 sky130_fd_sc_hd__nor2_1 _07028_ (.A(_01629_),
    .B(_01630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01631_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07029_ (.A(\sa_inst.sak._00_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01632_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07030_ (.A(_01632_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01633_));
 sky130_fd_sc_hd__nand2_1 _07031_ (.A(_01615_),
    .B(_01633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01634_));
 sky130_fd_sc_hd__xnor2_1 _07032_ (.A(_01631_),
    .B(_01634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01635_));
 sky130_fd_sc_hd__xnor2_1 _07033_ (.A(_01622_),
    .B(_01635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01636_));
 sky130_fd_sc_hd__xnor2_1 _07034_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._01_ ),
    .B(_01636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01637_));
 sky130_fd_sc_hd__mux2_1 _07035_ (.A0(_01624_),
    .A1(_01637_),
    .S(_01626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01638_));
 sky130_fd_sc_hd__clkbuf_1 _07036_ (.A(_01638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[2] ));
 sky130_fd_sc_hd__buf_2 _07037_ (.A(_01264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01639_));
 sky130_fd_sc_hd__and2_1 _07038_ (.A(_01622_),
    .B(_01635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01640_));
 sky130_fd_sc_hd__clkbuf_2 _07039_ (.A(\sa_inst._06_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01641_));
 sky130_fd_sc_hd__nand2_1 _07040_ (.A(_01614_),
    .B(_01641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01642_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07041_ (.A(\sa_inst.sak._00_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01643_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07042_ (.A(_01643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01644_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07043_ (.A(\sa_inst._06_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01645_));
 sky130_fd_sc_hd__a22oi_1 _07044_ (.A1(_01619_),
    .A2(_01645_),
    .B1(_01633_),
    .B2(_01618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01646_));
 sky130_fd_sc_hd__and3_1 _07045_ (.A(_01645_),
    .B(_01633_),
    .C(_01621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01647_));
 sky130_fd_sc_hd__o2bb2a_1 _07046_ (.A1_N(_01615_),
    .A2_N(_01644_),
    .B1(_01646_),
    .B2(_01647_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01648_));
 sky130_fd_sc_hd__and4bb_1 _07047_ (.A_N(_01646_),
    .B_N(_01647_),
    .C(\sa_inst._06_[4] ),
    .D(_01644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01649_));
 sky130_fd_sc_hd__nor2_1 _07048_ (.A(_01648_),
    .B(_01649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01650_));
 sky130_fd_sc_hd__xnor2_1 _07049_ (.A(_01642_),
    .B(_01650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01651_));
 sky130_fd_sc_hd__o21ba_1 _07050_ (.A1(_01630_),
    .A2(_01634_),
    .B1_N(_01629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01652_));
 sky130_fd_sc_hd__xnor2_1 _07051_ (.A(_01651_),
    .B(_01652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01653_));
 sky130_fd_sc_hd__and2_1 _07052_ (.A(_01640_),
    .B(_01653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01654_));
 sky130_fd_sc_hd__nor2_1 _07053_ (.A(_01640_),
    .B(_01653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01655_));
 sky130_fd_sc_hd__or2_1 _07054_ (.A(_01654_),
    .B(_01655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01656_));
 sky130_fd_sc_hd__xnor2_1 _07055_ (.A(_01639_),
    .B(_01656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01657_));
 sky130_fd_sc_hd__mux2_1 _07056_ (.A0(_01637_),
    .A1(_01657_),
    .S(_01626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01658_));
 sky130_fd_sc_hd__clkbuf_1 _07057_ (.A(_01658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[3] ));
 sky130_fd_sc_hd__and2b_1 _07058_ (.A_N(_01652_),
    .B(_01651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01659_));
 sky130_fd_sc_hd__or3_1 _07059_ (.A(_01642_),
    .B(_01648_),
    .C(_01649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01660_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07060_ (.A(\sa_inst._06_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01661_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07061_ (.A(_01661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01662_));
 sky130_fd_sc_hd__a22oi_1 _07062_ (.A1(_01619_),
    .A2(_01641_),
    .B1(_01662_),
    .B2(_01613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01663_));
 sky130_fd_sc_hd__and4_1 _07063_ (.A(_01613_),
    .B(_01619_),
    .C(\sa_inst._06_[7] ),
    .D(_01661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01664_));
 sky130_fd_sc_hd__nor2_1 _07064_ (.A(_01663_),
    .B(_01664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01665_));
 sky130_fd_sc_hd__a22oi_1 _07065_ (.A1(_01645_),
    .A2(_01632_),
    .B1(_01643_),
    .B2(\sa_inst._06_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01666_));
 sky130_fd_sc_hd__and4_1 _07066_ (.A(\sa_inst._06_[5] ),
    .B(\sa_inst._06_[6] ),
    .C(_01632_),
    .D(\sa_inst.sak._00_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01667_));
 sky130_fd_sc_hd__nor2_1 _07067_ (.A(_01666_),
    .B(_01667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01668_));
 sky130_fd_sc_hd__nand2_1 _07068_ (.A(\sa_inst._06_[4] ),
    .B(\sa_inst.sak._00_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01669_));
 sky130_fd_sc_hd__xnor2_1 _07069_ (.A(_01668_),
    .B(_01669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01670_));
 sky130_fd_sc_hd__xnor2_1 _07070_ (.A(_01665_),
    .B(_01670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01671_));
 sky130_fd_sc_hd__and2_1 _07071_ (.A(_01660_),
    .B(_01671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01672_));
 sky130_fd_sc_hd__nor2_1 _07072_ (.A(_01660_),
    .B(_01671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01673_));
 sky130_fd_sc_hd__nor2_1 _07073_ (.A(_01672_),
    .B(_01673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01674_));
 sky130_fd_sc_hd__or2_1 _07074_ (.A(_01647_),
    .B(_01649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01675_));
 sky130_fd_sc_hd__xor2_1 _07075_ (.A(_01674_),
    .B(_01675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01676_));
 sky130_fd_sc_hd__o21ai_2 _07076_ (.A1(_01659_),
    .A2(_01654_),
    .B1(_01676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01677_));
 sky130_fd_sc_hd__or3_1 _07077_ (.A(_01659_),
    .B(_01654_),
    .C(_01676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01678_));
 sky130_fd_sc_hd__nand2_1 _07078_ (.A(_01677_),
    .B(_01678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01679_));
 sky130_fd_sc_hd__xnor2_1 _07079_ (.A(_01639_),
    .B(_01679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01680_));
 sky130_fd_sc_hd__mux2_1 _07080_ (.A0(_01657_),
    .A1(_01680_),
    .S(_01626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01681_));
 sky130_fd_sc_hd__clkbuf_1 _07081_ (.A(_01681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[4] ));
 sky130_fd_sc_hd__and2_1 _07082_ (.A(_01665_),
    .B(_01670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01682_));
 sky130_fd_sc_hd__a22oi_1 _07083_ (.A1(\sa_inst.sak._00_[5] ),
    .A2(\sa_inst._06_[8] ),
    .B1(\sa_inst._06_[9] ),
    .B2(_01613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01683_));
 sky130_fd_sc_hd__and4_1 _07084_ (.A(\sa_inst.sak._00_[4] ),
    .B(\sa_inst.sak._00_[5] ),
    .C(\sa_inst._06_[8] ),
    .D(\sa_inst._06_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01684_));
 sky130_fd_sc_hd__o2bb2a_1 _07085_ (.A1_N(_01632_),
    .A2_N(\sa_inst._06_[7] ),
    .B1(_01683_),
    .B2(_01684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01685_));
 sky130_fd_sc_hd__and4bb_1 _07086_ (.A_N(_01683_),
    .B_N(_01684_),
    .C(_01632_),
    .D(\sa_inst._06_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01686_));
 sky130_fd_sc_hd__nor2_1 _07087_ (.A(_01685_),
    .B(_01686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01687_));
 sky130_fd_sc_hd__xnor2_1 _07088_ (.A(_01664_),
    .B(_01687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01688_));
 sky130_fd_sc_hd__a22oi_2 _07089_ (.A1(_01645_),
    .A2(_01643_),
    .B1(\sa_inst.sak._00_[8] ),
    .B2(_01618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01689_));
 sky130_fd_sc_hd__and4_1 _07090_ (.A(\sa_inst._06_[5] ),
    .B(\sa_inst._06_[6] ),
    .C(_01643_),
    .D(\sa_inst.sak._00_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01690_));
 sky130_fd_sc_hd__nand2_1 _07091_ (.A(\sa_inst._06_[4] ),
    .B(\sa_inst.sak._00_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01691_));
 sky130_fd_sc_hd__o21a_1 _07092_ (.A1(_01689_),
    .A2(_01690_),
    .B1(_01691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01692_));
 sky130_fd_sc_hd__nor3_2 _07093_ (.A(_01689_),
    .B(_01690_),
    .C(_01691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01693_));
 sky130_fd_sc_hd__nor2_1 _07094_ (.A(_01692_),
    .B(_01693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01694_));
 sky130_fd_sc_hd__xnor2_1 _07095_ (.A(_01688_),
    .B(_01694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01695_));
 sky130_fd_sc_hd__xnor2_1 _07096_ (.A(_01682_),
    .B(_01695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01696_));
 sky130_fd_sc_hd__o21ba_1 _07097_ (.A1(_01666_),
    .A2(_01669_),
    .B1_N(_01667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01697_));
 sky130_fd_sc_hd__xnor2_1 _07098_ (.A(_01696_),
    .B(_01697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01698_));
 sky130_fd_sc_hd__a21oi_1 _07099_ (.A1(_01674_),
    .A2(_01675_),
    .B1(_01673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01699_));
 sky130_fd_sc_hd__xnor2_1 _07100_ (.A(_01698_),
    .B(_01699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01700_));
 sky130_fd_sc_hd__xnor2_1 _07101_ (.A(_01677_),
    .B(_01700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01701_));
 sky130_fd_sc_hd__xnor2_1 _07102_ (.A(_01639_),
    .B(_01701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01702_));
 sky130_fd_sc_hd__clkbuf_2 _07103_ (.A(_01625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _07104_ (.A0(_01680_),
    .A1(_01702_),
    .S(_01703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01704_));
 sky130_fd_sc_hd__clkbuf_1 _07105_ (.A(_01704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[5] ));
 sky130_fd_sc_hd__nand2_1 _07106_ (.A(_01664_),
    .B(_01687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01705_));
 sky130_fd_sc_hd__or3_1 _07107_ (.A(_01688_),
    .B(_01692_),
    .C(_01693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01706_));
 sky130_fd_sc_hd__clkbuf_2 _07108_ (.A(\sa_inst._06_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01707_));
 sky130_fd_sc_hd__a22oi_1 _07109_ (.A1(\sa_inst.sak._00_[6] ),
    .A2(_01661_),
    .B1(_01707_),
    .B2(\sa_inst.sak._00_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01708_));
 sky130_fd_sc_hd__and4_1 _07110_ (.A(\sa_inst.sak._00_[5] ),
    .B(\sa_inst.sak._00_[6] ),
    .C(_01661_),
    .D(\sa_inst._06_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01709_));
 sky130_fd_sc_hd__nor2_1 _07111_ (.A(_01708_),
    .B(_01709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01710_));
 sky130_fd_sc_hd__nand2_1 _07112_ (.A(\sa_inst._06_[7] ),
    .B(\sa_inst.sak._00_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01711_));
 sky130_fd_sc_hd__xnor2_1 _07113_ (.A(_01710_),
    .B(_01711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01712_));
 sky130_fd_sc_hd__or2_1 _07114_ (.A(_01684_),
    .B(_01686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01713_));
 sky130_fd_sc_hd__xor2_1 _07115_ (.A(_01712_),
    .B(_01713_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01714_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07116_ (.A(\sa_inst.sak._00_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01715_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07117_ (.A(\sa_inst.sak._00_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01716_));
 sky130_fd_sc_hd__a22oi_1 _07118_ (.A1(_01628_),
    .A2(_01715_),
    .B1(_01716_),
    .B2(_01618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01717_));
 sky130_fd_sc_hd__and4_1 _07119_ (.A(_01618_),
    .B(_01645_),
    .C(\sa_inst.sak._00_[8] ),
    .D(\sa_inst.sak._00_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01718_));
 sky130_fd_sc_hd__nor2_1 _07120_ (.A(_01717_),
    .B(_01718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01719_));
 sky130_fd_sc_hd__xnor2_1 _07121_ (.A(_01714_),
    .B(_01719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01720_));
 sky130_fd_sc_hd__a21o_1 _07122_ (.A1(_01705_),
    .A2(_01706_),
    .B1(_01720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01721_));
 sky130_fd_sc_hd__nand3_1 _07123_ (.A(_01705_),
    .B(_01706_),
    .C(_01720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01722_));
 sky130_fd_sc_hd__o211ai_2 _07124_ (.A1(_01690_),
    .A2(_01693_),
    .B1(_01721_),
    .C1(_01722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01723_));
 sky130_fd_sc_hd__a211o_1 _07125_ (.A1(_01721_),
    .A2(_01722_),
    .B1(_01690_),
    .C1(_01693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01724_));
 sky130_fd_sc_hd__nand2_1 _07126_ (.A(_01682_),
    .B(_01695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01725_));
 sky130_fd_sc_hd__o21ai_1 _07127_ (.A1(_01696_),
    .A2(_01697_),
    .B1(_01725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01726_));
 sky130_fd_sc_hd__and3_1 _07128_ (.A(_01723_),
    .B(_01724_),
    .C(_01726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01727_));
 sky130_fd_sc_hd__a21oi_1 _07129_ (.A1(_01723_),
    .A2(_01724_),
    .B1(_01726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01728_));
 sky130_fd_sc_hd__or2_1 _07130_ (.A(_01727_),
    .B(_01728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01729_));
 sky130_fd_sc_hd__nor2_1 _07131_ (.A(_01698_),
    .B(_01699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01730_));
 sky130_fd_sc_hd__o21bai_1 _07132_ (.A1(_01677_),
    .A2(_01700_),
    .B1_N(_01730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01731_));
 sky130_fd_sc_hd__and2b_1 _07133_ (.A_N(_01729_),
    .B(_01731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01732_));
 sky130_fd_sc_hd__and2b_1 _07134_ (.A_N(_01731_),
    .B(_01729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01733_));
 sky130_fd_sc_hd__or2_1 _07135_ (.A(_01732_),
    .B(_01733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01734_));
 sky130_fd_sc_hd__xnor2_1 _07136_ (.A(_01639_),
    .B(_01734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01735_));
 sky130_fd_sc_hd__mux2_1 _07137_ (.A0(_01702_),
    .A1(_01735_),
    .S(_01703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01736_));
 sky130_fd_sc_hd__clkbuf_1 _07138_ (.A(_01736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[6] ));
 sky130_fd_sc_hd__nand2_1 _07139_ (.A(_01628_),
    .B(_01716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01737_));
 sky130_fd_sc_hd__a22oi_1 _07140_ (.A1(_01644_),
    .A2(_01662_),
    .B1(_01707_),
    .B2(_01633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01738_));
 sky130_fd_sc_hd__and4_1 _07141_ (.A(_01633_),
    .B(_01643_),
    .C(_01661_),
    .D(_01707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01739_));
 sky130_fd_sc_hd__nor2_1 _07142_ (.A(_01738_),
    .B(_01739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01740_));
 sky130_fd_sc_hd__nand2_1 _07143_ (.A(_01641_),
    .B(_01715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01741_));
 sky130_fd_sc_hd__xnor2_2 _07144_ (.A(_01740_),
    .B(_01741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01742_));
 sky130_fd_sc_hd__o21ba_1 _07145_ (.A1(_01708_),
    .A2(_01711_),
    .B1_N(_01709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01743_));
 sky130_fd_sc_hd__xnor2_2 _07146_ (.A(_01742_),
    .B(_01743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01744_));
 sky130_fd_sc_hd__xor2_2 _07147_ (.A(_01737_),
    .B(_01744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01745_));
 sky130_fd_sc_hd__a22o_1 _07148_ (.A1(_01712_),
    .A2(_01713_),
    .B1(_01714_),
    .B2(_01719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01746_));
 sky130_fd_sc_hd__xnor2_2 _07149_ (.A(_01745_),
    .B(_01746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01747_));
 sky130_fd_sc_hd__xnor2_2 _07150_ (.A(_01718_),
    .B(_01747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01748_));
 sky130_fd_sc_hd__nand2_1 _07151_ (.A(_01721_),
    .B(_01723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01749_));
 sky130_fd_sc_hd__xnor2_2 _07152_ (.A(_01748_),
    .B(_01749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01750_));
 sky130_fd_sc_hd__or3_1 _07153_ (.A(_01727_),
    .B(_01732_),
    .C(_01750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01751_));
 sky130_fd_sc_hd__o21ai_2 _07154_ (.A1(_01727_),
    .A2(_01732_),
    .B1(_01750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01752_));
 sky130_fd_sc_hd__nand2_1 _07155_ (.A(_01751_),
    .B(_01752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01753_));
 sky130_fd_sc_hd__xnor2_1 _07156_ (.A(_01639_),
    .B(_01753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01754_));
 sky130_fd_sc_hd__mux2_1 _07157_ (.A0(_01735_),
    .A1(_01754_),
    .S(_01703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01755_));
 sky130_fd_sc_hd__clkbuf_1 _07158_ (.A(_01755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[7] ));
 sky130_fd_sc_hd__a21o_1 _07159_ (.A1(_01721_),
    .A2(_01723_),
    .B1(_01748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01756_));
 sky130_fd_sc_hd__clkbuf_1 _07160_ (.A(_01707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01757_));
 sky130_fd_sc_hd__and2_1 _07161_ (.A(_01662_),
    .B(_01715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01758_));
 sky130_fd_sc_hd__a21oi_1 _07162_ (.A1(_01644_),
    .A2(_01757_),
    .B1(_01758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01759_));
 sky130_fd_sc_hd__and3_1 _07163_ (.A(_01644_),
    .B(_01707_),
    .C(_01758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01760_));
 sky130_fd_sc_hd__nor2_1 _07164_ (.A(_01759_),
    .B(_01760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01761_));
 sky130_fd_sc_hd__nand2_1 _07165_ (.A(_01641_),
    .B(_01716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01762_));
 sky130_fd_sc_hd__xnor2_1 _07166_ (.A(_01761_),
    .B(_01762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01763_));
 sky130_fd_sc_hd__o21ba_1 _07167_ (.A1(_01738_),
    .A2(_01741_),
    .B1_N(_01739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01764_));
 sky130_fd_sc_hd__inv_2 _07168_ (.A(_01764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01765_));
 sky130_fd_sc_hd__xnor2_1 _07169_ (.A(_01763_),
    .B(_01765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01766_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07170_ (.A(_01716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01767_));
 sky130_fd_sc_hd__and2b_1 _07171_ (.A_N(_01743_),
    .B(_01742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01768_));
 sky130_fd_sc_hd__a31oi_2 _07172_ (.A1(_01628_),
    .A2(_01767_),
    .A3(_01744_),
    .B1(_01768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01769_));
 sky130_fd_sc_hd__nor2_1 _07173_ (.A(_01766_),
    .B(_01769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01770_));
 sky130_fd_sc_hd__and2_1 _07174_ (.A(_01766_),
    .B(_01769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01771_));
 sky130_fd_sc_hd__and2b_1 _07175_ (.A_N(_01745_),
    .B(_01746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01772_));
 sky130_fd_sc_hd__a21oi_1 _07176_ (.A1(_01718_),
    .A2(_01747_),
    .B1(_01772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01773_));
 sky130_fd_sc_hd__or3_1 _07177_ (.A(_01770_),
    .B(_01771_),
    .C(_01773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01774_));
 sky130_fd_sc_hd__nor2_1 _07178_ (.A(_01770_),
    .B(_01771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01775_));
 sky130_fd_sc_hd__or2b_1 _07179_ (.A(_01775_),
    .B_N(_01773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01776_));
 sky130_fd_sc_hd__nand2_1 _07180_ (.A(_01774_),
    .B(_01776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01777_));
 sky130_fd_sc_hd__a21oi_1 _07181_ (.A1(_01756_),
    .A2(_01752_),
    .B1(_01777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01778_));
 sky130_fd_sc_hd__and3_1 _07182_ (.A(_01756_),
    .B(_01752_),
    .C(_01777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01779_));
 sky130_fd_sc_hd__nor2_1 _07183_ (.A(_01778_),
    .B(_01779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01780_));
 sky130_fd_sc_hd__xor2_1 _07184_ (.A(_01264_),
    .B(_01780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01781_));
 sky130_fd_sc_hd__mux2_1 _07185_ (.A0(_01754_),
    .A1(_01781_),
    .S(_01703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01782_));
 sky130_fd_sc_hd__clkbuf_1 _07186_ (.A(_01782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[8] ));
 sky130_fd_sc_hd__a21o_1 _07187_ (.A1(_01756_),
    .A2(_01752_),
    .B1(_01777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01783_));
 sky130_fd_sc_hd__a31o_1 _07188_ (.A1(_01641_),
    .A2(_01767_),
    .A3(_01761_),
    .B1(_01760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01784_));
 sky130_fd_sc_hd__a22oi_1 _07189_ (.A1(_01715_),
    .A2(_01757_),
    .B1(_01767_),
    .B2(_01662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01785_));
 sky130_fd_sc_hd__and4_1 _07190_ (.A(_01662_),
    .B(_01715_),
    .C(_01757_),
    .D(_01716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01786_));
 sky130_fd_sc_hd__nor2_1 _07191_ (.A(_01785_),
    .B(_01786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01787_));
 sky130_fd_sc_hd__xnor2_1 _07192_ (.A(_01784_),
    .B(_01787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01788_));
 sky130_fd_sc_hd__a21oi_1 _07193_ (.A1(_01763_),
    .A2(_01765_),
    .B1(_01770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01789_));
 sky130_fd_sc_hd__xnor2_1 _07194_ (.A(_01788_),
    .B(_01789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01790_));
 sky130_fd_sc_hd__a21oi_1 _07195_ (.A1(_01774_),
    .A2(_01783_),
    .B1(_01790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01791_));
 sky130_fd_sc_hd__and3_1 _07196_ (.A(_01774_),
    .B(_01783_),
    .C(_01790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01792_));
 sky130_fd_sc_hd__or2_1 _07197_ (.A(_01791_),
    .B(_01792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01793_));
 sky130_fd_sc_hd__xnor2_1 _07198_ (.A(_01264_),
    .B(_01793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01794_));
 sky130_fd_sc_hd__mux2_1 _07199_ (.A0(_01781_),
    .A1(_01794_),
    .S(_01703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01795_));
 sky130_fd_sc_hd__clkbuf_1 _07200_ (.A(_01795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[9] ));
 sky130_fd_sc_hd__inv_2 _07201_ (.A(_01788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01796_));
 sky130_fd_sc_hd__a21o_1 _07202_ (.A1(_01770_),
    .A2(_01796_),
    .B1(_01791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01797_));
 sky130_fd_sc_hd__and3b_1 _07203_ (.A_N(_01758_),
    .B(_01767_),
    .C(_01757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01798_));
 sky130_fd_sc_hd__and2_1 _07204_ (.A(_01784_),
    .B(_01787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01799_));
 sky130_fd_sc_hd__and3_1 _07205_ (.A(_01763_),
    .B(_01765_),
    .C(_01796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01800_));
 sky130_fd_sc_hd__nor2_1 _07206_ (.A(_01799_),
    .B(_01800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01801_));
 sky130_fd_sc_hd__xnor2_1 _07207_ (.A(_01798_),
    .B(_01801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01802_));
 sky130_fd_sc_hd__xnor2_1 _07208_ (.A(_01797_),
    .B(_01802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01803_));
 sky130_fd_sc_hd__xnor2_1 _07209_ (.A(_01264_),
    .B(_01803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01804_));
 sky130_fd_sc_hd__mux2_1 _07210_ (.A0(_01794_),
    .A1(_01804_),
    .S(_01625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01805_));
 sky130_fd_sc_hd__clkbuf_1 _07211_ (.A(_01805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[10] ));
 sky130_fd_sc_hd__a22o_1 _07212_ (.A1(_01798_),
    .A2(_01800_),
    .B1(_01802_),
    .B2(_01797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01806_));
 sky130_fd_sc_hd__o211a_1 _07213_ (.A1(_01758_),
    .A2(_01799_),
    .B1(_01757_),
    .C1(_01767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01807_));
 sky130_fd_sc_hd__xnor2_1 _07214_ (.A(_01263_),
    .B(_01807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01808_));
 sky130_fd_sc_hd__xnor2_1 _07215_ (.A(_01806_),
    .B(_01808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01809_));
 sky130_fd_sc_hd__mux2_1 _07216_ (.A0(_01804_),
    .A1(_01809_),
    .S(_01625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01810_));
 sky130_fd_sc_hd__clkbuf_1 _07217_ (.A(_01810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[11] ));
 sky130_fd_sc_hd__mux2_1 _07218_ (.A0(_01809_),
    .A1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._01_ ),
    .S(_01625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01811_));
 sky130_fd_sc_hd__clkbuf_1 _07219_ (.A(_01811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[12] ));
 sky130_fd_sc_hd__xor2_1 _07220_ (.A(\sa_inst._07_[10] ),
    .B(\sa_inst.sak._08_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01812_));
 sky130_fd_sc_hd__clkbuf_2 _07221_ (.A(_01812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01813_));
 sky130_fd_sc_hd__clkbuf_2 _07222_ (.A(_01813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._01_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07223_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._00_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01814_));
 sky130_fd_sc_hd__clkbuf_4 _07224_ (.A(_01814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01815_));
 sky130_fd_sc_hd__inv_2 _07225_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01816_));
 sky130_fd_sc_hd__clkbuf_2 _07226_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01817_));
 sky130_fd_sc_hd__mux2_1 _07227_ (.A0(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ),
    .A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[1] ),
    .S(_01817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01818_));
 sky130_fd_sc_hd__and2b_1 _07228_ (.A_N(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._22_ ),
    .B(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01819_));
 sky130_fd_sc_hd__mux4_2 _07229_ (.A0(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .A2(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .A3(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .S0(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ),
    .S1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01820_));
 sky130_fd_sc_hd__clkbuf_2 _07230_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01821_));
 sky130_fd_sc_hd__nor2_1 _07231_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._22_ ),
    .B(_01821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01822_));
 sky130_fd_sc_hd__a32o_2 _07232_ (.A1(_01816_),
    .A2(_01818_),
    .A3(_01819_),
    .B1(_01820_),
    .B2(_01822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01823_));
 sky130_fd_sc_hd__xor2_4 _07233_ (.A(_01815_),
    .B(_01823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01824_));
 sky130_fd_sc_hd__clkbuf_1 _07234_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01825_));
 sky130_fd_sc_hd__clkbuf_4 _07235_ (.A(_01825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01826_));
 sky130_fd_sc_hd__nand2_1 _07236_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[0] ),
    .B(_01826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01827_));
 sky130_fd_sc_hd__xnor2_1 _07237_ (.A(_01824_),
    .B(_01827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[0] ));
 sky130_fd_sc_hd__clkbuf_4 _07238_ (.A(_01825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01828_));
 sky130_fd_sc_hd__clkbuf_4 _07239_ (.A(_01828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01829_));
 sky130_fd_sc_hd__inv_2 _07240_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._22_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01830_));
 sky130_fd_sc_hd__clkbuf_2 _07241_ (.A(_01830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _07242_ (.A0(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .S(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _07243_ (.A0(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .S(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01833_));
 sky130_fd_sc_hd__mux2_1 _07244_ (.A0(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ),
    .A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[2] ),
    .S(_01817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01834_));
 sky130_fd_sc_hd__clkbuf_2 _07245_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01835_));
 sky130_fd_sc_hd__and2b_1 _07246_ (.A_N(_01835_),
    .B(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01836_));
 sky130_fd_sc_hd__buf_2 _07247_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01837_));
 sky130_fd_sc_hd__mux4_2 _07248_ (.A0(_01832_),
    .A1(_01833_),
    .A2(_01834_),
    .A3(_01836_),
    .S0(_01837_),
    .S1(_01821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01838_));
 sky130_fd_sc_hd__nand4_4 _07249_ (.A(_01831_),
    .B(_01815_),
    .C(_01823_),
    .D(_01838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01839_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07250_ (.A(_01839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01840_));
 sky130_fd_sc_hd__clkbuf_2 _07251_ (.A(_01831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01841_));
 sky130_fd_sc_hd__a22o_1 _07252_ (.A1(_01815_),
    .A2(_01823_),
    .B1(_01838_),
    .B2(_01841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01842_));
 sky130_fd_sc_hd__and3_1 _07253_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[1] ),
    .B(_01840_),
    .C(_01842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01843_));
 sky130_fd_sc_hd__a21oi_1 _07254_ (.A1(_01840_),
    .A2(_01842_),
    .B1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01844_));
 sky130_fd_sc_hd__or2_1 _07255_ (.A(_01843_),
    .B(_01844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01845_));
 sky130_fd_sc_hd__nand2_1 _07256_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[0] ),
    .B(_01824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01846_));
 sky130_fd_sc_hd__or2_1 _07257_ (.A(_01845_),
    .B(_01846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01847_));
 sky130_fd_sc_hd__nand2_1 _07258_ (.A(_01845_),
    .B(_01846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01848_));
 sky130_fd_sc_hd__inv_2 _07259_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01849_));
 sky130_fd_sc_hd__clkbuf_2 _07260_ (.A(_01849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01850_));
 sky130_fd_sc_hd__and3_1 _07261_ (.A(_01850_),
    .B(_01840_),
    .C(_01842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01851_));
 sky130_fd_sc_hd__a31o_1 _07262_ (.A1(_01829_),
    .A2(_01847_),
    .A3(_01848_),
    .B1(_01851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[1] ));
 sky130_fd_sc_hd__o21ba_1 _07263_ (.A1(_01844_),
    .A2(_01846_),
    .B1_N(_01843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01852_));
 sky130_fd_sc_hd__clkbuf_2 _07264_ (.A(_01817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01853_));
 sky130_fd_sc_hd__mux4_2 _07265_ (.A0(_01814_),
    .A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .A2(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .A3(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .S0(_01837_),
    .S1(_01853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01854_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07266_ (.A(_01816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _07267_ (.A0(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ),
    .S(_01853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01856_));
 sky130_fd_sc_hd__clkbuf_2 _07268_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01857_));
 sky130_fd_sc_hd__and3b_1 _07269_ (.A_N(_01853_),
    .B(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[1] ),
    .C(_01857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01858_));
 sky130_fd_sc_hd__a21o_1 _07270_ (.A1(_01855_),
    .A2(_01856_),
    .B1(_01858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01859_));
 sky130_fd_sc_hd__a22oi_4 _07271_ (.A1(_01822_),
    .A2(_01854_),
    .B1(_01859_),
    .B2(_01819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01860_));
 sky130_fd_sc_hd__xor2_2 _07272_ (.A(_01839_),
    .B(_01860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01861_));
 sky130_fd_sc_hd__nor2_1 _07273_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[2] ),
    .B(_01861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01862_));
 sky130_fd_sc_hd__clkbuf_1 _07274_ (.A(_01861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01863_));
 sky130_fd_sc_hd__and2_1 _07275_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[2] ),
    .B(_01863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01864_));
 sky130_fd_sc_hd__or3_1 _07276_ (.A(_01852_),
    .B(_01862_),
    .C(_01864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01865_));
 sky130_fd_sc_hd__o21ai_1 _07277_ (.A1(_01862_),
    .A2(_01864_),
    .B1(_01852_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01866_));
 sky130_fd_sc_hd__clkbuf_2 _07278_ (.A(_01850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01867_));
 sky130_fd_sc_hd__and2_1 _07279_ (.A(_01867_),
    .B(_01863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01868_));
 sky130_fd_sc_hd__a31o_1 _07280_ (.A1(_01829_),
    .A2(_01865_),
    .A3(_01866_),
    .B1(_01868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[2] ));
 sky130_fd_sc_hd__mux4_2 _07281_ (.A0(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._00_ ),
    .A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .A2(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .A3(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .S0(_01837_),
    .S1(_01853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01869_));
 sky130_fd_sc_hd__mux4_1 _07282_ (.A0(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[2] ),
    .A2(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ),
    .A3(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[0] ),
    .S0(_01837_),
    .S1(_01853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01870_));
 sky130_fd_sc_hd__a22o_1 _07283_ (.A1(_01822_),
    .A2(_01869_),
    .B1(_01870_),
    .B2(_01819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01871_));
 sky130_fd_sc_hd__nor3b_1 _07284_ (.A(_01839_),
    .B(_01860_),
    .C_N(_01871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01872_));
 sky130_fd_sc_hd__buf_2 _07285_ (.A(_01872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01873_));
 sky130_fd_sc_hd__clkbuf_2 _07286_ (.A(_01873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01874_));
 sky130_fd_sc_hd__o21ba_1 _07287_ (.A1(_01840_),
    .A2(_01860_),
    .B1_N(_01871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01875_));
 sky130_fd_sc_hd__nor2_1 _07288_ (.A(_01874_),
    .B(_01875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01876_));
 sky130_fd_sc_hd__nor2_1 _07289_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[3] ),
    .B(_01876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01877_));
 sky130_fd_sc_hd__or3b_1 _07290_ (.A(_01873_),
    .B(_01875_),
    .C_N(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01878_));
 sky130_fd_sc_hd__or2b_1 _07291_ (.A(_01877_),
    .B_N(_01878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01879_));
 sky130_fd_sc_hd__nand2_1 _07292_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[2] ),
    .B(_01863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01880_));
 sky130_fd_sc_hd__o21ai_1 _07293_ (.A1(_01852_),
    .A2(_01862_),
    .B1(_01880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01881_));
 sky130_fd_sc_hd__xnor2_1 _07294_ (.A(_01879_),
    .B(_01881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01882_));
 sky130_fd_sc_hd__buf_2 _07295_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _07296_ (.A0(_01876_),
    .A1(_01882_),
    .S(_01883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01884_));
 sky130_fd_sc_hd__clkbuf_1 _07297_ (.A(_01884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[3] ));
 sky130_fd_sc_hd__mux2_1 _07298_ (.A0(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .S(_01817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01885_));
 sky130_fd_sc_hd__mux2_1 _07299_ (.A0(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .S(_01817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01886_));
 sky130_fd_sc_hd__mux4_1 _07300_ (.A0(_01814_),
    .A1(_01885_),
    .A2(_01886_),
    .A3(_01818_),
    .S0(_01857_),
    .S1(_01821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01887_));
 sky130_fd_sc_hd__and2_1 _07301_ (.A(_01841_),
    .B(_01887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01888_));
 sky130_fd_sc_hd__xor2_4 _07302_ (.A(_01873_),
    .B(_01888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01889_));
 sky130_fd_sc_hd__xnor2_1 _07303_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[4] ),
    .B(_01889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01890_));
 sky130_fd_sc_hd__o211a_1 _07304_ (.A1(_01852_),
    .A2(_01862_),
    .B1(_01880_),
    .C1(_01878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01891_));
 sky130_fd_sc_hd__or3_1 _07305_ (.A(_01877_),
    .B(_01890_),
    .C(_01891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01892_));
 sky130_fd_sc_hd__o21ai_1 _07306_ (.A1(_01877_),
    .A2(_01891_),
    .B1(_01890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01893_));
 sky130_fd_sc_hd__and2_1 _07307_ (.A(_01867_),
    .B(_01889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01894_));
 sky130_fd_sc_hd__a31o_1 _07308_ (.A1(_01829_),
    .A2(_01892_),
    .A3(_01893_),
    .B1(_01894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[4] ));
 sky130_fd_sc_hd__mux4_1 _07309_ (.A0(_01814_),
    .A1(_01832_),
    .A2(_01833_),
    .A3(_01834_),
    .S0(_01857_),
    .S1(_01821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01895_));
 sky130_fd_sc_hd__a22o_1 _07310_ (.A1(_01873_),
    .A2(_01888_),
    .B1(_01895_),
    .B2(_01841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01896_));
 sky130_fd_sc_hd__and3_1 _07311_ (.A(_01831_),
    .B(_01887_),
    .C(_01895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01897_));
 sky130_fd_sc_hd__nand2_1 _07312_ (.A(_01874_),
    .B(_01897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01898_));
 sky130_fd_sc_hd__and2_1 _07313_ (.A(_01896_),
    .B(_01898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01899_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07314_ (.A(_01899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01900_));
 sky130_fd_sc_hd__nand2_1 _07315_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[5] ),
    .B(_01899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01901_));
 sky130_fd_sc_hd__clkinv_2 _07316_ (.A(_01901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01902_));
 sky130_fd_sc_hd__nor2_1 _07317_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[5] ),
    .B(_01900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01903_));
 sky130_fd_sc_hd__or2_1 _07318_ (.A(_01902_),
    .B(_01903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01904_));
 sky130_fd_sc_hd__and2_1 _07319_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[4] ),
    .B(_01889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01905_));
 sky130_fd_sc_hd__inv_2 _07320_ (.A(_01905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01906_));
 sky130_fd_sc_hd__and2_1 _07321_ (.A(_01906_),
    .B(_01892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01907_));
 sky130_fd_sc_hd__xor2_1 _07322_ (.A(_01904_),
    .B(_01907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01908_));
 sky130_fd_sc_hd__mux2_1 _07323_ (.A0(_01900_),
    .A1(_01908_),
    .S(_01883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01909_));
 sky130_fd_sc_hd__clkbuf_1 _07324_ (.A(_01909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[5] ));
 sky130_fd_sc_hd__buf_2 _07325_ (.A(_01849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01910_));
 sky130_fd_sc_hd__buf_2 _07326_ (.A(_01910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01911_));
 sky130_fd_sc_hd__clkbuf_2 _07327_ (.A(_01821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01912_));
 sky130_fd_sc_hd__mux2_1 _07328_ (.A0(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._00_ ),
    .A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .S(_01835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01913_));
 sky130_fd_sc_hd__nor2_1 _07329_ (.A(_01857_),
    .B(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._00_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01914_));
 sky130_fd_sc_hd__o21ba_1 _07330_ (.A1(_01855_),
    .A2(_01913_),
    .B1_N(_01914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01915_));
 sky130_fd_sc_hd__inv_2 _07331_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01916_));
 sky130_fd_sc_hd__mux4_1 _07332_ (.A0(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .A2(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .A3(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ),
    .S0(_01835_),
    .S1(_01837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01917_));
 sky130_fd_sc_hd__or2_1 _07333_ (.A(_01916_),
    .B(_01917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01918_));
 sky130_fd_sc_hd__o211a_1 _07334_ (.A1(_01912_),
    .A2(_01915_),
    .B1(_01918_),
    .C1(_01831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01919_));
 sky130_fd_sc_hd__xnor2_2 _07335_ (.A(_01898_),
    .B(_01919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01920_));
 sky130_fd_sc_hd__clkbuf_2 _07336_ (.A(_01920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01921_));
 sky130_fd_sc_hd__xnor2_1 _07337_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[6] ),
    .B(_01920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01922_));
 sky130_fd_sc_hd__a311o_1 _07338_ (.A1(_01906_),
    .A2(_01892_),
    .A3(_01901_),
    .B1(_01903_),
    .C1(_01922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01923_));
 sky130_fd_sc_hd__clkbuf_4 _07339_ (.A(_01849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01924_));
 sky130_fd_sc_hd__o211a_1 _07340_ (.A1(_01903_),
    .A2(_01907_),
    .B1(_01922_),
    .C1(_01901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01925_));
 sky130_fd_sc_hd__nor2_1 _07341_ (.A(_01924_),
    .B(_01925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01926_));
 sky130_fd_sc_hd__a22o_1 _07342_ (.A1(_01911_),
    .A2(_01921_),
    .B1(_01923_),
    .B2(_01926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[6] ));
 sky130_fd_sc_hd__clkbuf_2 _07343_ (.A(_01828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01927_));
 sky130_fd_sc_hd__mux2_1 _07344_ (.A0(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._00_ ),
    .A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .S(_01835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01928_));
 sky130_fd_sc_hd__o21ba_1 _07345_ (.A1(_01855_),
    .A2(_01928_),
    .B1_N(_01914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01929_));
 sky130_fd_sc_hd__mux4_1 _07346_ (.A0(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .A2(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .A3(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ),
    .S0(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .S1(_01835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01930_));
 sky130_fd_sc_hd__or2_1 _07347_ (.A(_01916_),
    .B(_01930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01931_));
 sky130_fd_sc_hd__o211a_1 _07348_ (.A1(_01912_),
    .A2(_01929_),
    .B1(_01931_),
    .C1(_01831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01932_));
 sky130_fd_sc_hd__and3_1 _07349_ (.A(_01897_),
    .B(_01919_),
    .C(_01932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01933_));
 sky130_fd_sc_hd__nand2_2 _07350_ (.A(_01874_),
    .B(_01933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01934_));
 sky130_fd_sc_hd__a31o_1 _07351_ (.A1(_01874_),
    .A2(_01897_),
    .A3(_01919_),
    .B1(_01932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01935_));
 sky130_fd_sc_hd__and2_2 _07352_ (.A(_01934_),
    .B(_01935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01936_));
 sky130_fd_sc_hd__nor2_1 _07353_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[7] ),
    .B(_01936_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01937_));
 sky130_fd_sc_hd__and3_1 _07354_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[7] ),
    .B(_01934_),
    .C(_01935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01938_));
 sky130_fd_sc_hd__or2_1 _07355_ (.A(_01937_),
    .B(_01938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01939_));
 sky130_fd_sc_hd__and2_1 _07356_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[6] ),
    .B(_01921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01940_));
 sky130_fd_sc_hd__or2b_1 _07357_ (.A(_01940_),
    .B_N(_01923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01941_));
 sky130_fd_sc_hd__xnor2_1 _07358_ (.A(_01939_),
    .B(_01941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01942_));
 sky130_fd_sc_hd__and3_1 _07359_ (.A(_01910_),
    .B(_01934_),
    .C(_01935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01943_));
 sky130_fd_sc_hd__a21o_1 _07360_ (.A1(_01927_),
    .A2(_01942_),
    .B1(_01943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[7] ));
 sky130_fd_sc_hd__or2_1 _07361_ (.A(_01916_),
    .B(_01820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01944_));
 sky130_fd_sc_hd__o21a_1 _07362_ (.A1(_01912_),
    .A2(_01814_),
    .B1(_01830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01945_));
 sky130_fd_sc_hd__and2_2 _07363_ (.A(_01944_),
    .B(_01945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01946_));
 sky130_fd_sc_hd__xnor2_4 _07364_ (.A(_01934_),
    .B(_01946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01947_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07365_ (.A(_01947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01948_));
 sky130_fd_sc_hd__xnor2_1 _07366_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[8] ),
    .B(_01947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01949_));
 sky130_fd_sc_hd__nor2_1 _07367_ (.A(_01940_),
    .B(_01938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01950_));
 sky130_fd_sc_hd__a21o_1 _07368_ (.A1(_01923_),
    .A2(_01950_),
    .B1(_01937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01951_));
 sky130_fd_sc_hd__or2_1 _07369_ (.A(_01949_),
    .B(_01951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01952_));
 sky130_fd_sc_hd__a21oi_1 _07370_ (.A1(_01949_),
    .A2(_01951_),
    .B1(_01924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01953_));
 sky130_fd_sc_hd__a22o_1 _07371_ (.A1(_01911_),
    .A2(_01948_),
    .B1(_01952_),
    .B2(_01953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[8] ));
 sky130_fd_sc_hd__mux2_1 _07372_ (.A0(_01832_),
    .A1(_01833_),
    .S(_01857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01954_));
 sky130_fd_sc_hd__o21a_1 _07373_ (.A1(_01916_),
    .A2(_01954_),
    .B1(_01945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01955_));
 sky130_fd_sc_hd__and2_1 _07374_ (.A(_01944_),
    .B(_01955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01956_));
 sky130_fd_sc_hd__nand3_2 _07375_ (.A(_01872_),
    .B(_01933_),
    .C(_01956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01957_));
 sky130_fd_sc_hd__clkbuf_2 _07376_ (.A(_01957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01958_));
 sky130_fd_sc_hd__a31o_1 _07377_ (.A1(_01874_),
    .A2(_01933_),
    .A3(_01946_),
    .B1(_01955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01959_));
 sky130_fd_sc_hd__and2_1 _07378_ (.A(_01958_),
    .B(_01959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01960_));
 sky130_fd_sc_hd__and3_1 _07379_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[9] ),
    .B(_01958_),
    .C(_01959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01961_));
 sky130_fd_sc_hd__a21oi_1 _07380_ (.A1(_01958_),
    .A2(_01959_),
    .B1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01962_));
 sky130_fd_sc_hd__or2_1 _07381_ (.A(_01961_),
    .B(_01962_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01963_));
 sky130_fd_sc_hd__a21bo_1 _07382_ (.A1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[8] ),
    .A2(_01948_),
    .B1_N(_01952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01964_));
 sky130_fd_sc_hd__xnor2_1 _07383_ (.A(_01963_),
    .B(_01964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01965_));
 sky130_fd_sc_hd__mux2_1 _07384_ (.A0(_01960_),
    .A1(_01965_),
    .S(_01883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01966_));
 sky130_fd_sc_hd__clkbuf_1 _07385_ (.A(_01966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[9] ));
 sky130_fd_sc_hd__o21ai_2 _07386_ (.A1(_01912_),
    .A2(_01815_),
    .B1(_01841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01967_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07387_ (.A(_01916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01968_));
 sky130_fd_sc_hd__nor2_1 _07388_ (.A(_01968_),
    .B(_01854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01969_));
 sky130_fd_sc_hd__or2_2 _07389_ (.A(_01967_),
    .B(_01969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01970_));
 sky130_fd_sc_hd__xor2_2 _07390_ (.A(_01957_),
    .B(_01970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01971_));
 sky130_fd_sc_hd__xnor2_1 _07391_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[10] ),
    .B(_01971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01972_));
 sky130_fd_sc_hd__a21oi_1 _07392_ (.A1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[8] ),
    .A2(_01947_),
    .B1(_01961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01973_));
 sky130_fd_sc_hd__a21o_1 _07393_ (.A1(_01952_),
    .A2(_01973_),
    .B1(_01962_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01974_));
 sky130_fd_sc_hd__xor2_1 _07394_ (.A(_01972_),
    .B(_01974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01975_));
 sky130_fd_sc_hd__clkbuf_2 _07395_ (.A(_01971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01976_));
 sky130_fd_sc_hd__and2_1 _07396_ (.A(_01910_),
    .B(_01976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01977_));
 sky130_fd_sc_hd__a21o_1 _07397_ (.A1(_01927_),
    .A2(_01975_),
    .B1(_01977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[10] ));
 sky130_fd_sc_hd__buf_2 _07398_ (.A(_01825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01978_));
 sky130_fd_sc_hd__buf_2 _07399_ (.A(_01978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01979_));
 sky130_fd_sc_hd__nor2_2 _07400_ (.A(_01968_),
    .B(_01869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01980_));
 sky130_fd_sc_hd__or3_1 _07401_ (.A(_01957_),
    .B(_01970_),
    .C(_01980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01981_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07402_ (.A(_01981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01982_));
 sky130_fd_sc_hd__o22ai_4 _07403_ (.A1(_01958_),
    .A2(_01970_),
    .B1(_01980_),
    .B2(_01967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01983_));
 sky130_fd_sc_hd__and3_1 _07404_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[11] ),
    .B(_01982_),
    .C(_01983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01984_));
 sky130_fd_sc_hd__a21oi_1 _07405_ (.A1(_01982_),
    .A2(_01983_),
    .B1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01985_));
 sky130_fd_sc_hd__or2_1 _07406_ (.A(_01984_),
    .B(_01985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01986_));
 sky130_fd_sc_hd__o2bb2ai_1 _07407_ (.A1_N(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[10] ),
    .A2_N(_01976_),
    .B1(_01972_),
    .B2(_01974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01987_));
 sky130_fd_sc_hd__xnor2_1 _07408_ (.A(_01986_),
    .B(_01987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01988_));
 sky130_fd_sc_hd__and3_1 _07409_ (.A(_01850_),
    .B(_01982_),
    .C(_01983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01989_));
 sky130_fd_sc_hd__a21o_1 _07410_ (.A1(_01979_),
    .A2(_01988_),
    .B1(_01989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[11] ));
 sky130_fd_sc_hd__clkbuf_2 _07411_ (.A(_01826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01990_));
 sky130_fd_sc_hd__a21o_1 _07412_ (.A1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[10] ),
    .A2(_01976_),
    .B1(_01984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01991_));
 sky130_fd_sc_hd__or2b_1 _07413_ (.A(_01985_),
    .B_N(_01991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01992_));
 sky130_fd_sc_hd__or3_1 _07414_ (.A(_01972_),
    .B(_01984_),
    .C(_01985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01993_));
 sky130_fd_sc_hd__or3_1 _07415_ (.A(_01962_),
    .B(_01973_),
    .C(_01993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01994_));
 sky130_fd_sc_hd__or2_1 _07416_ (.A(_01949_),
    .B(_01963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01995_));
 sky130_fd_sc_hd__a2111o_1 _07417_ (.A1(_01923_),
    .A2(_01950_),
    .B1(_01993_),
    .C1(_01995_),
    .D1(_01937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01996_));
 sky130_fd_sc_hd__o21ba_1 _07418_ (.A1(_01855_),
    .A2(_01885_),
    .B1_N(_01914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01997_));
 sky130_fd_sc_hd__o31a_1 _07419_ (.A1(_01957_),
    .A2(_01969_),
    .A3(_01980_),
    .B1(_01945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01998_));
 sky130_fd_sc_hd__clkbuf_2 _07420_ (.A(_01998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01999_));
 sky130_fd_sc_hd__o21a_1 _07421_ (.A1(_01968_),
    .A2(_01997_),
    .B1(_01999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02000_));
 sky130_fd_sc_hd__clkbuf_2 _07422_ (.A(_02000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02001_));
 sky130_fd_sc_hd__xnor2_1 _07423_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[12] ),
    .B(_02001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02002_));
 sky130_fd_sc_hd__a31o_1 _07424_ (.A1(_01992_),
    .A2(_01994_),
    .A3(_01996_),
    .B1(_02002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02003_));
 sky130_fd_sc_hd__nand4_1 _07425_ (.A(_02002_),
    .B(_01992_),
    .C(_01994_),
    .D(_01996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02004_));
 sky130_fd_sc_hd__and2_1 _07426_ (.A(_01867_),
    .B(_02001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02005_));
 sky130_fd_sc_hd__a31o_1 _07427_ (.A1(_01990_),
    .A2(_02003_),
    .A3(_02004_),
    .B1(_02005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[12] ));
 sky130_fd_sc_hd__nor2_1 _07428_ (.A(_01855_),
    .B(_01832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02006_));
 sky130_fd_sc_hd__o21ai_2 _07429_ (.A1(_01914_),
    .A2(_02006_),
    .B1(_01912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02007_));
 sky130_fd_sc_hd__and3_1 _07430_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[13] ),
    .B(_01999_),
    .C(_02007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02008_));
 sky130_fd_sc_hd__a21oi_1 _07431_ (.A1(_01999_),
    .A2(_02007_),
    .B1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02009_));
 sky130_fd_sc_hd__or2_1 _07432_ (.A(_02008_),
    .B(_02009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02010_));
 sky130_fd_sc_hd__a21bo_1 _07433_ (.A1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[12] ),
    .A2(_02001_),
    .B1_N(_02003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02011_));
 sky130_fd_sc_hd__xnor2_1 _07434_ (.A(_02010_),
    .B(_02011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02012_));
 sky130_fd_sc_hd__nand2_1 _07435_ (.A(_01999_),
    .B(_02007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02013_));
 sky130_fd_sc_hd__nor2_1 _07436_ (.A(_01978_),
    .B(_02013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02014_));
 sky130_fd_sc_hd__a21o_1 _07437_ (.A1(_01979_),
    .A2(_02012_),
    .B1(_02014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[13] ));
 sky130_fd_sc_hd__nor2_1 _07438_ (.A(_02008_),
    .B(_02011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02015_));
 sky130_fd_sc_hd__o21a_2 _07439_ (.A1(_01968_),
    .A2(_01915_),
    .B1(_01999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02016_));
 sky130_fd_sc_hd__xnor2_2 _07440_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[14] ),
    .B(_02016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02017_));
 sky130_fd_sc_hd__o21ai_1 _07441_ (.A1(_02009_),
    .A2(_02015_),
    .B1(_02017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02018_));
 sky130_fd_sc_hd__or2_1 _07442_ (.A(_02009_),
    .B(_02017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02019_));
 sky130_fd_sc_hd__or2_1 _07443_ (.A(_02015_),
    .B(_02019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02020_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07444_ (.A(_02016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02021_));
 sky130_fd_sc_hd__and2_1 _07445_ (.A(_01867_),
    .B(_02021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02022_));
 sky130_fd_sc_hd__a31o_1 _07446_ (.A1(_01990_),
    .A2(_02018_),
    .A3(_02020_),
    .B1(_02022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[14] ));
 sky130_fd_sc_hd__nand2_1 _07447_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[14] ),
    .B(_02021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02023_));
 sky130_fd_sc_hd__o21a_1 _07448_ (.A1(_01968_),
    .A2(_01929_),
    .B1(_01998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02024_));
 sky130_fd_sc_hd__and2_1 _07449_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[15] ),
    .B(_02024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02025_));
 sky130_fd_sc_hd__clkbuf_2 _07450_ (.A(_02024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02026_));
 sky130_fd_sc_hd__nor2_1 _07451_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[15] ),
    .B(_02026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02027_));
 sky130_fd_sc_hd__or2_2 _07452_ (.A(_02025_),
    .B(_02027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02028_));
 sky130_fd_sc_hd__a21o_1 _07453_ (.A1(_02023_),
    .A2(_02020_),
    .B1(_02028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02029_));
 sky130_fd_sc_hd__nand3_1 _07454_ (.A(_02023_),
    .B(_02020_),
    .C(_02028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02030_));
 sky130_fd_sc_hd__and2_1 _07455_ (.A(_01867_),
    .B(_02026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02031_));
 sky130_fd_sc_hd__a31o_1 _07456_ (.A1(_01990_),
    .A2(_02029_),
    .A3(_02030_),
    .B1(_02031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[15] ));
 sky130_fd_sc_hd__a21oi_1 _07457_ (.A1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[12] ),
    .A2(_02001_),
    .B1(_02008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02032_));
 sky130_fd_sc_hd__a21oi_1 _07458_ (.A1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[14] ),
    .A2(_02021_),
    .B1(_02025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02033_));
 sky130_fd_sc_hd__o32a_1 _07459_ (.A1(_02032_),
    .A2(_02019_),
    .A3(_02028_),
    .B1(_02033_),
    .B2(_02027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02034_));
 sky130_fd_sc_hd__o41ai_4 _07460_ (.A1(_02003_),
    .A2(_02010_),
    .A3(_02017_),
    .A4(_02028_),
    .B1(_02034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02035_));
 sky130_fd_sc_hd__and3_1 _07461_ (.A(_01841_),
    .B(_01815_),
    .C(_01981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02036_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07462_ (.A(_02036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02037_));
 sky130_fd_sc_hd__clkbuf_2 _07463_ (.A(_02037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02038_));
 sky130_fd_sc_hd__xnor2_1 _07464_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[16] ),
    .B(_02038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02039_));
 sky130_fd_sc_hd__xnor2_1 _07465_ (.A(_02035_),
    .B(_02039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02040_));
 sky130_fd_sc_hd__buf_2 _07466_ (.A(_02037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02041_));
 sky130_fd_sc_hd__buf_2 _07467_ (.A(_02041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02042_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07468_ (.A(_02042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02043_));
 sky130_fd_sc_hd__clkbuf_2 _07469_ (.A(_02043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02044_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07470_ (.A(_02044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02045_));
 sky130_fd_sc_hd__clkbuf_2 _07471_ (.A(_02045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02046_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07472_ (.A(_02046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02047_));
 sky130_fd_sc_hd__and2_1 _07473_ (.A(_01849_),
    .B(_02047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02048_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07474_ (.A(_02048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02049_));
 sky130_fd_sc_hd__buf_2 _07475_ (.A(_02049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02050_));
 sky130_fd_sc_hd__a21o_1 _07476_ (.A1(_01979_),
    .A2(_02040_),
    .B1(_02050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[16] ));
 sky130_fd_sc_hd__and2b_1 _07477_ (.A_N(_02039_),
    .B(_02035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02051_));
 sky130_fd_sc_hd__a21oi_1 _07478_ (.A1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[16] ),
    .A2(_02046_),
    .B1(_02051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02052_));
 sky130_fd_sc_hd__clkbuf_2 _07479_ (.A(_02037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02053_));
 sky130_fd_sc_hd__nand2_1 _07480_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[17] ),
    .B(_02053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02054_));
 sky130_fd_sc_hd__clkbuf_2 _07481_ (.A(_02036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02055_));
 sky130_fd_sc_hd__or2_1 _07482_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[17] ),
    .B(_02055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02056_));
 sky130_fd_sc_hd__nand2_1 _07483_ (.A(_02054_),
    .B(_02056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02057_));
 sky130_fd_sc_hd__or2_1 _07484_ (.A(_02052_),
    .B(_02057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02058_));
 sky130_fd_sc_hd__nand2_1 _07485_ (.A(_02052_),
    .B(_02057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02059_));
 sky130_fd_sc_hd__buf_2 _07486_ (.A(_02049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02060_));
 sky130_fd_sc_hd__a31o_1 _07487_ (.A1(_01990_),
    .A2(_02058_),
    .A3(_02059_),
    .B1(_02060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[17] ));
 sky130_fd_sc_hd__or2b_1 _07488_ (.A(_02052_),
    .B_N(_02056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02061_));
 sky130_fd_sc_hd__nand2_1 _07489_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[18] ),
    .B(_02038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02062_));
 sky130_fd_sc_hd__or2_1 _07490_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[18] ),
    .B(_02041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02063_));
 sky130_fd_sc_hd__nand2_1 _07491_ (.A(_02062_),
    .B(_02063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02064_));
 sky130_fd_sc_hd__a21o_1 _07492_ (.A1(_02054_),
    .A2(_02061_),
    .B1(_02064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02065_));
 sky130_fd_sc_hd__nand3_1 _07493_ (.A(_02054_),
    .B(_02061_),
    .C(_02064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02066_));
 sky130_fd_sc_hd__a31o_1 _07494_ (.A1(_01990_),
    .A2(_02065_),
    .A3(_02066_),
    .B1(_02060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[18] ));
 sky130_fd_sc_hd__clkbuf_2 _07495_ (.A(_01826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02067_));
 sky130_fd_sc_hd__xnor2_1 _07496_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[19] ),
    .B(_02038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02068_));
 sky130_fd_sc_hd__a21o_1 _07497_ (.A1(_02062_),
    .A2(_02065_),
    .B1(_02068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02069_));
 sky130_fd_sc_hd__nand3_1 _07498_ (.A(_02062_),
    .B(_02065_),
    .C(_02068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02070_));
 sky130_fd_sc_hd__clkbuf_2 _07499_ (.A(_02049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02071_));
 sky130_fd_sc_hd__a31o_1 _07500_ (.A1(_02067_),
    .A2(_02069_),
    .A3(_02070_),
    .B1(_02071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[19] ));
 sky130_fd_sc_hd__nand2_1 _07501_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[20] ),
    .B(_02038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02072_));
 sky130_fd_sc_hd__or2_1 _07502_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[20] ),
    .B(_02041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02073_));
 sky130_fd_sc_hd__nand2_1 _07503_ (.A(_02072_),
    .B(_02073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02074_));
 sky130_fd_sc_hd__or4_1 _07504_ (.A(_02039_),
    .B(_02057_),
    .C(_02064_),
    .D(_02068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02075_));
 sky130_fd_sc_hd__inv_2 _07505_ (.A(_02075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02076_));
 sky130_fd_sc_hd__buf_2 _07506_ (.A(_02043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02077_));
 sky130_fd_sc_hd__o41a_1 _07507_ (.A1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[16] ),
    .A2(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[17] ),
    .A3(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[18] ),
    .A4(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[19] ),
    .B1(_02077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02078_));
 sky130_fd_sc_hd__a21oi_1 _07508_ (.A1(_02035_),
    .A2(_02076_),
    .B1(_02078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02079_));
 sky130_fd_sc_hd__or2_1 _07509_ (.A(_02074_),
    .B(_02079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02080_));
 sky130_fd_sc_hd__nand2_1 _07510_ (.A(_02074_),
    .B(_02079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02081_));
 sky130_fd_sc_hd__a31o_1 _07511_ (.A1(_02067_),
    .A2(_02080_),
    .A3(_02081_),
    .B1(_02071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[20] ));
 sky130_fd_sc_hd__o21a_1 _07512_ (.A1(_02074_),
    .A2(_02079_),
    .B1(_02072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02082_));
 sky130_fd_sc_hd__nand2_1 _07513_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[21] ),
    .B(_02038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02083_));
 sky130_fd_sc_hd__or2_1 _07514_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[21] ),
    .B(_02041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02084_));
 sky130_fd_sc_hd__nand2_1 _07515_ (.A(_02083_),
    .B(_02084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02085_));
 sky130_fd_sc_hd__or2_1 _07516_ (.A(_02082_),
    .B(_02085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02086_));
 sky130_fd_sc_hd__nand2_1 _07517_ (.A(_02082_),
    .B(_02085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02087_));
 sky130_fd_sc_hd__a31o_1 _07518_ (.A1(_02067_),
    .A2(_02086_),
    .A3(_02087_),
    .B1(_02071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[21] ));
 sky130_fd_sc_hd__or2b_1 _07519_ (.A(_02082_),
    .B_N(_02084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02088_));
 sky130_fd_sc_hd__and2_1 _07520_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[22] ),
    .B(_02055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02089_));
 sky130_fd_sc_hd__nor2_1 _07521_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[22] ),
    .B(_02053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02090_));
 sky130_fd_sc_hd__or2_1 _07522_ (.A(_02089_),
    .B(_02090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02091_));
 sky130_fd_sc_hd__a21oi_1 _07523_ (.A1(_02083_),
    .A2(_02088_),
    .B1(_02091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02092_));
 sky130_fd_sc_hd__clkbuf_4 _07524_ (.A(_01850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02093_));
 sky130_fd_sc_hd__a31o_1 _07525_ (.A1(_02083_),
    .A2(_02088_),
    .A3(_02091_),
    .B1(_02093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02094_));
 sky130_fd_sc_hd__clkbuf_2 _07526_ (.A(_02048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02095_));
 sky130_fd_sc_hd__o21bai_1 _07527_ (.A1(_02092_),
    .A2(_02094_),
    .B1_N(_02095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[22] ));
 sky130_fd_sc_hd__xor2_1 _07528_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[23] ),
    .B(_02042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02096_));
 sky130_fd_sc_hd__o21ai_1 _07529_ (.A1(_02089_),
    .A2(_02092_),
    .B1(_02096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02097_));
 sky130_fd_sc_hd__or3_1 _07530_ (.A(_02089_),
    .B(_02092_),
    .C(_02096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02098_));
 sky130_fd_sc_hd__a31o_1 _07531_ (.A1(_02067_),
    .A2(_02097_),
    .A3(_02098_),
    .B1(_02071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[23] ));
 sky130_fd_sc_hd__or4b_1 _07532_ (.A(_02074_),
    .B(_02085_),
    .C(_02091_),
    .D_N(_02096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02099_));
 sky130_fd_sc_hd__nor2_1 _07533_ (.A(_02075_),
    .B(_02099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02100_));
 sky130_fd_sc_hd__o41a_1 _07534_ (.A1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[20] ),
    .A2(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[21] ),
    .A3(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[22] ),
    .A4(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[23] ),
    .B1(_02077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02101_));
 sky130_fd_sc_hd__a211o_2 _07535_ (.A1(_02035_),
    .A2(_02100_),
    .B1(_02101_),
    .C1(_02078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02102_));
 sky130_fd_sc_hd__xor2_2 _07536_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[24] ),
    .B(_02077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02103_));
 sky130_fd_sc_hd__nand2_1 _07537_ (.A(_02102_),
    .B(_02103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02104_));
 sky130_fd_sc_hd__o21a_1 _07538_ (.A1(_02102_),
    .A2(_02103_),
    .B1(_01828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02105_));
 sky130_fd_sc_hd__a21o_1 _07539_ (.A1(_02104_),
    .A2(_02105_),
    .B1(_02050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[24] ));
 sky130_fd_sc_hd__xor2_1 _07540_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[25] ),
    .B(_02077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02106_));
 sky130_fd_sc_hd__clkbuf_4 _07541_ (.A(_02047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02107_));
 sky130_fd_sc_hd__a22o_1 _07542_ (.A1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[24] ),
    .A2(_02107_),
    .B1(_02102_),
    .B2(_02103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02108_));
 sky130_fd_sc_hd__xor2_1 _07543_ (.A(_02106_),
    .B(_02108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02109_));
 sky130_fd_sc_hd__a21o_1 _07544_ (.A1(_01979_),
    .A2(_02109_),
    .B1(_02050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[25] ));
 sky130_fd_sc_hd__clkbuf_2 _07545_ (.A(_02045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02110_));
 sky130_fd_sc_hd__o21ai_1 _07546_ (.A1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[24] ),
    .A2(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[25] ),
    .B1(_02110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02111_));
 sky130_fd_sc_hd__and2_1 _07547_ (.A(_02103_),
    .B(_02106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02112_));
 sky130_fd_sc_hd__nand2_1 _07548_ (.A(_02102_),
    .B(_02112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02113_));
 sky130_fd_sc_hd__nand2_1 _07549_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[26] ),
    .B(_02044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02114_));
 sky130_fd_sc_hd__or2_1 _07550_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[26] ),
    .B(_02043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02115_));
 sky130_fd_sc_hd__nand2_1 _07551_ (.A(_02114_),
    .B(_02115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02116_));
 sky130_fd_sc_hd__a21o_1 _07552_ (.A1(_02111_),
    .A2(_02113_),
    .B1(_02116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02117_));
 sky130_fd_sc_hd__nand3_1 _07553_ (.A(_02116_),
    .B(_02111_),
    .C(_02113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02118_));
 sky130_fd_sc_hd__a31o_1 _07554_ (.A1(_02067_),
    .A2(_02117_),
    .A3(_02118_),
    .B1(_02071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[26] ));
 sky130_fd_sc_hd__xnor2_1 _07555_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[27] ),
    .B(_02044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02119_));
 sky130_fd_sc_hd__nand2_1 _07556_ (.A(_02114_),
    .B(_02117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02120_));
 sky130_fd_sc_hd__xnor2_1 _07557_ (.A(_02119_),
    .B(_02120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02121_));
 sky130_fd_sc_hd__a21o_1 _07558_ (.A1(_01979_),
    .A2(_02121_),
    .B1(_02050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[27] ));
 sky130_fd_sc_hd__nor2_1 _07559_ (.A(_02116_),
    .B(_02119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02122_));
 sky130_fd_sc_hd__clkbuf_2 _07560_ (.A(_02043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02123_));
 sky130_fd_sc_hd__clkbuf_2 _07561_ (.A(_02123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02124_));
 sky130_fd_sc_hd__o41a_1 _07562_ (.A1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[24] ),
    .A2(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[25] ),
    .A3(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[26] ),
    .A4(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[27] ),
    .B1(_02124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02125_));
 sky130_fd_sc_hd__a31oi_2 _07563_ (.A1(_02102_),
    .A2(_02112_),
    .A3(_02122_),
    .B1(_02125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02126_));
 sky130_fd_sc_hd__and2_1 _07564_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[28] ),
    .B(_02124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02127_));
 sky130_fd_sc_hd__nor2_1 _07565_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[28] ),
    .B(_02124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02128_));
 sky130_fd_sc_hd__or2_1 _07566_ (.A(_02127_),
    .B(_02128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02129_));
 sky130_fd_sc_hd__nor2_1 _07567_ (.A(_02126_),
    .B(_02129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02130_));
 sky130_fd_sc_hd__a21o_1 _07568_ (.A1(_02126_),
    .A2(_02129_),
    .B1(_01924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02131_));
 sky130_fd_sc_hd__o21bai_1 _07569_ (.A1(_02130_),
    .A2(_02131_),
    .B1_N(_02095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[28] ));
 sky130_fd_sc_hd__buf_2 _07570_ (.A(_01826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02132_));
 sky130_fd_sc_hd__nand2_1 _07571_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[29] ),
    .B(_02046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02133_));
 sky130_fd_sc_hd__or2_1 _07572_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[29] ),
    .B(_02045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02134_));
 sky130_fd_sc_hd__o211ai_1 _07573_ (.A1(_02127_),
    .A2(_02130_),
    .B1(_02133_),
    .C1(_02134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02135_));
 sky130_fd_sc_hd__a211o_1 _07574_ (.A1(_02133_),
    .A2(_02134_),
    .B1(_02127_),
    .C1(_02130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02136_));
 sky130_fd_sc_hd__clkbuf_2 _07575_ (.A(_02048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02137_));
 sky130_fd_sc_hd__a31o_1 _07576_ (.A1(_02132_),
    .A2(_02135_),
    .A3(_02136_),
    .B1(_02137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[29] ));
 sky130_fd_sc_hd__o21ai_1 _07577_ (.A1(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[28] ),
    .A2(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[29] ),
    .B1(_02047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02138_));
 sky130_fd_sc_hd__or4bb_1 _07578_ (.A(_02126_),
    .B(_02129_),
    .C_N(_02133_),
    .D_N(_02134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02139_));
 sky130_fd_sc_hd__and2_1 _07579_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[30] ),
    .B(_02046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02140_));
 sky130_fd_sc_hd__nor2_1 _07580_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[30] ),
    .B(_02110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02141_));
 sky130_fd_sc_hd__or2_1 _07581_ (.A(_02140_),
    .B(_02141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02142_));
 sky130_fd_sc_hd__a21o_1 _07582_ (.A1(_02138_),
    .A2(_02139_),
    .B1(_02142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02143_));
 sky130_fd_sc_hd__nand3_1 _07583_ (.A(_02142_),
    .B(_02138_),
    .C(_02139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02144_));
 sky130_fd_sc_hd__a31o_1 _07584_ (.A1(_02132_),
    .A2(_02143_),
    .A3(_02144_),
    .B1(_02137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[30] ));
 sky130_fd_sc_hd__nand2_1 _07585_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[31] ),
    .B(_02107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02145_));
 sky130_fd_sc_hd__or2_1 _07586_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[31] ),
    .B(_02047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02146_));
 sky130_fd_sc_hd__a21oi_1 _07587_ (.A1(_02138_),
    .A2(_02139_),
    .B1(_02142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02147_));
 sky130_fd_sc_hd__a211o_1 _07588_ (.A1(_02145_),
    .A2(_02146_),
    .B1(_02140_),
    .C1(_02147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02148_));
 sky130_fd_sc_hd__o211ai_1 _07589_ (.A1(_02140_),
    .A2(_02147_),
    .B1(_02145_),
    .C1(_02146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02149_));
 sky130_fd_sc_hd__a31o_1 _07590_ (.A1(_02132_),
    .A2(_02148_),
    .A3(_02149_),
    .B1(_02137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[31] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07591_ (.A(\sa_inst._07_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02150_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07592_ (.A(\sa_inst.sak._08_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02151_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07593_ (.A(_02151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02152_));
 sky130_fd_sc_hd__nand2_1 _07594_ (.A(_02150_),
    .B(_02152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02153_));
 sky130_fd_sc_hd__xnor2_1 _07595_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._01_ ),
    .B(_02153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02154_));
 sky130_fd_sc_hd__clkbuf_2 _07596_ (.A(\sa_inst._07_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02155_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07597_ (.A(\sa_inst.sak._08_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02156_));
 sky130_fd_sc_hd__a22oi_1 _07598_ (.A1(_02152_),
    .A2(_02155_),
    .B1(_02156_),
    .B2(_02150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02157_));
 sky130_fd_sc_hd__and2_1 _07599_ (.A(\sa_inst._07_[5] ),
    .B(_02156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02158_));
 sky130_fd_sc_hd__and3_1 _07600_ (.A(_02150_),
    .B(_02152_),
    .C(_02158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02159_));
 sky130_fd_sc_hd__or2_1 _07601_ (.A(_02157_),
    .B(_02159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02160_));
 sky130_fd_sc_hd__xnor2_1 _07602_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._01_ ),
    .B(_02160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02161_));
 sky130_fd_sc_hd__xor2_4 _07603_ (.A(\sa_inst._07_[0] ),
    .B(\sa_inst.sak._08_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02162_));
 sky130_fd_sc_hd__clkbuf_2 _07604_ (.A(_02162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02163_));
 sky130_fd_sc_hd__mux2_1 _07605_ (.A0(_02154_),
    .A1(_02161_),
    .S(_02163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02164_));
 sky130_fd_sc_hd__clkbuf_1 _07606_ (.A(_02164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[1] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07607_ (.A(\sa_inst._07_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02165_));
 sky130_fd_sc_hd__and3_1 _07608_ (.A(_02151_),
    .B(_02165_),
    .C(_02158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02166_));
 sky130_fd_sc_hd__a21oi_1 _07609_ (.A1(_02152_),
    .A2(_02165_),
    .B1(_02158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02167_));
 sky130_fd_sc_hd__nor2_1 _07610_ (.A(_02166_),
    .B(_02167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02168_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07611_ (.A(\sa_inst.sak._08_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02169_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07612_ (.A(_02169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02170_));
 sky130_fd_sc_hd__nand2_1 _07613_ (.A(_02150_),
    .B(_02170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02171_));
 sky130_fd_sc_hd__xnor2_1 _07614_ (.A(_02168_),
    .B(_02171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02172_));
 sky130_fd_sc_hd__xnor2_1 _07615_ (.A(_02159_),
    .B(_02172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02173_));
 sky130_fd_sc_hd__xnor2_1 _07616_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._01_ ),
    .B(_02173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02174_));
 sky130_fd_sc_hd__mux2_1 _07617_ (.A0(_02161_),
    .A1(_02174_),
    .S(_02163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02175_));
 sky130_fd_sc_hd__clkbuf_1 _07618_ (.A(_02175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[2] ));
 sky130_fd_sc_hd__buf_2 _07619_ (.A(_01813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02176_));
 sky130_fd_sc_hd__and2_1 _07620_ (.A(_02159_),
    .B(_02172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02177_));
 sky130_fd_sc_hd__clkbuf_2 _07621_ (.A(\sa_inst._07_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02178_));
 sky130_fd_sc_hd__nand2_1 _07622_ (.A(_02152_),
    .B(_02178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02179_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07623_ (.A(\sa_inst.sak._08_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02180_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07624_ (.A(_02180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02181_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07625_ (.A(\sa_inst._07_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02182_));
 sky130_fd_sc_hd__a22oi_1 _07626_ (.A1(_02156_),
    .A2(_02182_),
    .B1(_02170_),
    .B2(_02155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02183_));
 sky130_fd_sc_hd__and3_1 _07627_ (.A(_02182_),
    .B(_02170_),
    .C(_02158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02184_));
 sky130_fd_sc_hd__o2bb2a_1 _07628_ (.A1_N(_02150_),
    .A2_N(_02181_),
    .B1(_02183_),
    .B2(_02184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02185_));
 sky130_fd_sc_hd__and4bb_1 _07629_ (.A_N(_02183_),
    .B_N(_02184_),
    .C(\sa_inst._07_[4] ),
    .D(_02181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02186_));
 sky130_fd_sc_hd__nor2_1 _07630_ (.A(_02185_),
    .B(_02186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02187_));
 sky130_fd_sc_hd__xnor2_1 _07631_ (.A(_02179_),
    .B(_02187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02188_));
 sky130_fd_sc_hd__o21ba_1 _07632_ (.A1(_02167_),
    .A2(_02171_),
    .B1_N(_02166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02189_));
 sky130_fd_sc_hd__xnor2_1 _07633_ (.A(_02188_),
    .B(_02189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02190_));
 sky130_fd_sc_hd__and2_1 _07634_ (.A(_02177_),
    .B(_02190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02191_));
 sky130_fd_sc_hd__nor2_1 _07635_ (.A(_02177_),
    .B(_02190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02192_));
 sky130_fd_sc_hd__or2_1 _07636_ (.A(_02191_),
    .B(_02192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02193_));
 sky130_fd_sc_hd__xnor2_1 _07637_ (.A(_02176_),
    .B(_02193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02194_));
 sky130_fd_sc_hd__mux2_1 _07638_ (.A0(_02174_),
    .A1(_02194_),
    .S(_02163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02195_));
 sky130_fd_sc_hd__clkbuf_1 _07639_ (.A(_02195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[3] ));
 sky130_fd_sc_hd__and2b_1 _07640_ (.A_N(_02189_),
    .B(_02188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02196_));
 sky130_fd_sc_hd__or3_1 _07641_ (.A(_02179_),
    .B(_02185_),
    .C(_02186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02197_));
 sky130_fd_sc_hd__clkbuf_1 _07642_ (.A(\sa_inst._07_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02198_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07643_ (.A(_02198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02199_));
 sky130_fd_sc_hd__a22oi_1 _07644_ (.A1(_02156_),
    .A2(_02178_),
    .B1(_02199_),
    .B2(_02151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02200_));
 sky130_fd_sc_hd__and4_1 _07645_ (.A(_02151_),
    .B(_02156_),
    .C(\sa_inst._07_[7] ),
    .D(_02198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02201_));
 sky130_fd_sc_hd__nor2_1 _07646_ (.A(_02200_),
    .B(_02201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02202_));
 sky130_fd_sc_hd__a22oi_1 _07647_ (.A1(_02182_),
    .A2(_02169_),
    .B1(_02180_),
    .B2(\sa_inst._07_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02203_));
 sky130_fd_sc_hd__and4_1 _07648_ (.A(\sa_inst._07_[5] ),
    .B(\sa_inst._07_[6] ),
    .C(_02169_),
    .D(\sa_inst.sak._08_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02204_));
 sky130_fd_sc_hd__nor2_1 _07649_ (.A(_02203_),
    .B(_02204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02205_));
 sky130_fd_sc_hd__nand2_1 _07650_ (.A(\sa_inst._07_[4] ),
    .B(\sa_inst.sak._08_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02206_));
 sky130_fd_sc_hd__xnor2_1 _07651_ (.A(_02205_),
    .B(_02206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02207_));
 sky130_fd_sc_hd__xnor2_1 _07652_ (.A(_02202_),
    .B(_02207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02208_));
 sky130_fd_sc_hd__and2_1 _07653_ (.A(_02197_),
    .B(_02208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02209_));
 sky130_fd_sc_hd__nor2_1 _07654_ (.A(_02197_),
    .B(_02208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02210_));
 sky130_fd_sc_hd__nor2_1 _07655_ (.A(_02209_),
    .B(_02210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02211_));
 sky130_fd_sc_hd__or2_1 _07656_ (.A(_02184_),
    .B(_02186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02212_));
 sky130_fd_sc_hd__xor2_1 _07657_ (.A(_02211_),
    .B(_02212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02213_));
 sky130_fd_sc_hd__o21ai_2 _07658_ (.A1(_02196_),
    .A2(_02191_),
    .B1(_02213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02214_));
 sky130_fd_sc_hd__or3_1 _07659_ (.A(_02196_),
    .B(_02191_),
    .C(_02213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02215_));
 sky130_fd_sc_hd__nand2_1 _07660_ (.A(_02214_),
    .B(_02215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02216_));
 sky130_fd_sc_hd__xnor2_1 _07661_ (.A(_02176_),
    .B(_02216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02217_));
 sky130_fd_sc_hd__mux2_1 _07662_ (.A0(_02194_),
    .A1(_02217_),
    .S(_02163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02218_));
 sky130_fd_sc_hd__clkbuf_1 _07663_ (.A(_02218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[4] ));
 sky130_fd_sc_hd__and2_1 _07664_ (.A(_02202_),
    .B(_02207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02219_));
 sky130_fd_sc_hd__a22oi_1 _07665_ (.A1(\sa_inst.sak._08_[5] ),
    .A2(\sa_inst._07_[8] ),
    .B1(\sa_inst._07_[9] ),
    .B2(_02151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02220_));
 sky130_fd_sc_hd__and4_1 _07666_ (.A(\sa_inst.sak._08_[4] ),
    .B(\sa_inst.sak._08_[5] ),
    .C(\sa_inst._07_[8] ),
    .D(\sa_inst._07_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02221_));
 sky130_fd_sc_hd__o2bb2a_1 _07667_ (.A1_N(_02169_),
    .A2_N(\sa_inst._07_[7] ),
    .B1(_02220_),
    .B2(_02221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02222_));
 sky130_fd_sc_hd__and4bb_1 _07668_ (.A_N(_02220_),
    .B_N(_02221_),
    .C(_02169_),
    .D(\sa_inst._07_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02223_));
 sky130_fd_sc_hd__nor2_1 _07669_ (.A(_02222_),
    .B(_02223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02224_));
 sky130_fd_sc_hd__xnor2_1 _07670_ (.A(_02201_),
    .B(_02224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02225_));
 sky130_fd_sc_hd__a22oi_2 _07671_ (.A1(_02182_),
    .A2(_02180_),
    .B1(\sa_inst.sak._08_[8] ),
    .B2(_02155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02226_));
 sky130_fd_sc_hd__and4_1 _07672_ (.A(\sa_inst._07_[5] ),
    .B(\sa_inst._07_[6] ),
    .C(_02180_),
    .D(\sa_inst.sak._08_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02227_));
 sky130_fd_sc_hd__nand2_1 _07673_ (.A(\sa_inst._07_[4] ),
    .B(\sa_inst.sak._08_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02228_));
 sky130_fd_sc_hd__o21a_1 _07674_ (.A1(_02226_),
    .A2(_02227_),
    .B1(_02228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02229_));
 sky130_fd_sc_hd__nor3_1 _07675_ (.A(_02226_),
    .B(_02227_),
    .C(_02228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02230_));
 sky130_fd_sc_hd__nor2_1 _07676_ (.A(_02229_),
    .B(_02230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02231_));
 sky130_fd_sc_hd__xnor2_1 _07677_ (.A(_02225_),
    .B(_02231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02232_));
 sky130_fd_sc_hd__xnor2_1 _07678_ (.A(_02219_),
    .B(_02232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02233_));
 sky130_fd_sc_hd__o21ba_1 _07679_ (.A1(_02203_),
    .A2(_02206_),
    .B1_N(_02204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02234_));
 sky130_fd_sc_hd__xnor2_1 _07680_ (.A(_02233_),
    .B(_02234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02235_));
 sky130_fd_sc_hd__a21oi_1 _07681_ (.A1(_02211_),
    .A2(_02212_),
    .B1(_02210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02236_));
 sky130_fd_sc_hd__xnor2_1 _07682_ (.A(_02235_),
    .B(_02236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02237_));
 sky130_fd_sc_hd__xnor2_1 _07683_ (.A(_02214_),
    .B(_02237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02238_));
 sky130_fd_sc_hd__xnor2_1 _07684_ (.A(_02176_),
    .B(_02238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02239_));
 sky130_fd_sc_hd__clkbuf_2 _07685_ (.A(_02162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02240_));
 sky130_fd_sc_hd__mux2_1 _07686_ (.A0(_02217_),
    .A1(_02239_),
    .S(_02240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02241_));
 sky130_fd_sc_hd__clkbuf_1 _07687_ (.A(_02241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[5] ));
 sky130_fd_sc_hd__nand2_1 _07688_ (.A(_02201_),
    .B(_02224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02242_));
 sky130_fd_sc_hd__or3_1 _07689_ (.A(_02225_),
    .B(_02229_),
    .C(_02230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02243_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07690_ (.A(\sa_inst._07_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02244_));
 sky130_fd_sc_hd__a22oi_1 _07691_ (.A1(\sa_inst.sak._08_[6] ),
    .A2(_02198_),
    .B1(_02244_),
    .B2(\sa_inst.sak._08_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02245_));
 sky130_fd_sc_hd__and4_1 _07692_ (.A(\sa_inst.sak._08_[5] ),
    .B(\sa_inst.sak._08_[6] ),
    .C(_02198_),
    .D(\sa_inst._07_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02246_));
 sky130_fd_sc_hd__nor2_1 _07693_ (.A(_02245_),
    .B(_02246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02247_));
 sky130_fd_sc_hd__nand2_1 _07694_ (.A(\sa_inst._07_[7] ),
    .B(\sa_inst.sak._08_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02248_));
 sky130_fd_sc_hd__xnor2_1 _07695_ (.A(_02247_),
    .B(_02248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02249_));
 sky130_fd_sc_hd__or2_1 _07696_ (.A(_02221_),
    .B(_02223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02250_));
 sky130_fd_sc_hd__xor2_1 _07697_ (.A(_02249_),
    .B(_02250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02251_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07698_ (.A(\sa_inst.sak._08_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02252_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07699_ (.A(\sa_inst.sak._08_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02253_));
 sky130_fd_sc_hd__a22oi_1 _07700_ (.A1(_02165_),
    .A2(_02252_),
    .B1(_02253_),
    .B2(_02155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02254_));
 sky130_fd_sc_hd__and4_1 _07701_ (.A(_02155_),
    .B(_02182_),
    .C(\sa_inst.sak._08_[8] ),
    .D(\sa_inst.sak._08_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02255_));
 sky130_fd_sc_hd__nor2_1 _07702_ (.A(_02254_),
    .B(_02255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02256_));
 sky130_fd_sc_hd__xnor2_1 _07703_ (.A(_02251_),
    .B(_02256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02257_));
 sky130_fd_sc_hd__a21o_1 _07704_ (.A1(_02242_),
    .A2(_02243_),
    .B1(_02257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02258_));
 sky130_fd_sc_hd__nand3_1 _07705_ (.A(_02242_),
    .B(_02243_),
    .C(_02257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02259_));
 sky130_fd_sc_hd__o211ai_2 _07706_ (.A1(_02227_),
    .A2(_02230_),
    .B1(_02258_),
    .C1(_02259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02260_));
 sky130_fd_sc_hd__a211o_1 _07707_ (.A1(_02258_),
    .A2(_02259_),
    .B1(_02227_),
    .C1(_02230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02261_));
 sky130_fd_sc_hd__nand2_1 _07708_ (.A(_02219_),
    .B(_02232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02262_));
 sky130_fd_sc_hd__o21ai_1 _07709_ (.A1(_02233_),
    .A2(_02234_),
    .B1(_02262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02263_));
 sky130_fd_sc_hd__and3_1 _07710_ (.A(_02260_),
    .B(_02261_),
    .C(_02263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02264_));
 sky130_fd_sc_hd__a21oi_1 _07711_ (.A1(_02260_),
    .A2(_02261_),
    .B1(_02263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02265_));
 sky130_fd_sc_hd__or2_1 _07712_ (.A(_02264_),
    .B(_02265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02266_));
 sky130_fd_sc_hd__nor2_1 _07713_ (.A(_02235_),
    .B(_02236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02267_));
 sky130_fd_sc_hd__o21bai_1 _07714_ (.A1(_02214_),
    .A2(_02237_),
    .B1_N(_02267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02268_));
 sky130_fd_sc_hd__and2b_1 _07715_ (.A_N(_02266_),
    .B(_02268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02269_));
 sky130_fd_sc_hd__and2b_1 _07716_ (.A_N(_02268_),
    .B(_02266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02270_));
 sky130_fd_sc_hd__or2_1 _07717_ (.A(_02269_),
    .B(_02270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02271_));
 sky130_fd_sc_hd__xnor2_1 _07718_ (.A(_02176_),
    .B(_02271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02272_));
 sky130_fd_sc_hd__mux2_1 _07719_ (.A0(_02239_),
    .A1(_02272_),
    .S(_02240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02273_));
 sky130_fd_sc_hd__clkbuf_1 _07720_ (.A(_02273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[6] ));
 sky130_fd_sc_hd__nand2_1 _07721_ (.A(_02165_),
    .B(_02253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02274_));
 sky130_fd_sc_hd__a22oi_1 _07722_ (.A1(_02181_),
    .A2(_02199_),
    .B1(_02244_),
    .B2(_02170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02275_));
 sky130_fd_sc_hd__and4_1 _07723_ (.A(_02170_),
    .B(_02180_),
    .C(_02198_),
    .D(_02244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02276_));
 sky130_fd_sc_hd__nor2_1 _07724_ (.A(_02275_),
    .B(_02276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02277_));
 sky130_fd_sc_hd__nand2_1 _07725_ (.A(_02178_),
    .B(_02252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02278_));
 sky130_fd_sc_hd__xnor2_1 _07726_ (.A(_02277_),
    .B(_02278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02279_));
 sky130_fd_sc_hd__o21ba_1 _07727_ (.A1(_02245_),
    .A2(_02248_),
    .B1_N(_02246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02280_));
 sky130_fd_sc_hd__xnor2_1 _07728_ (.A(_02279_),
    .B(_02280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02281_));
 sky130_fd_sc_hd__xor2_1 _07729_ (.A(_02274_),
    .B(_02281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02282_));
 sky130_fd_sc_hd__a22o_1 _07730_ (.A1(_02249_),
    .A2(_02250_),
    .B1(_02251_),
    .B2(_02256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02283_));
 sky130_fd_sc_hd__xnor2_1 _07731_ (.A(_02282_),
    .B(_02283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02284_));
 sky130_fd_sc_hd__xnor2_1 _07732_ (.A(_02255_),
    .B(_02284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02285_));
 sky130_fd_sc_hd__nand2_1 _07733_ (.A(_02258_),
    .B(_02260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02286_));
 sky130_fd_sc_hd__xnor2_1 _07734_ (.A(_02285_),
    .B(_02286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02287_));
 sky130_fd_sc_hd__or3_1 _07735_ (.A(_02264_),
    .B(_02269_),
    .C(_02287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02288_));
 sky130_fd_sc_hd__o21ai_2 _07736_ (.A1(_02264_),
    .A2(_02269_),
    .B1(_02287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02289_));
 sky130_fd_sc_hd__nand2_1 _07737_ (.A(_02288_),
    .B(_02289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02290_));
 sky130_fd_sc_hd__xnor2_1 _07738_ (.A(_02176_),
    .B(_02290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02291_));
 sky130_fd_sc_hd__mux2_1 _07739_ (.A0(_02272_),
    .A1(_02291_),
    .S(_02240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02292_));
 sky130_fd_sc_hd__clkbuf_1 _07740_ (.A(_02292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[7] ));
 sky130_fd_sc_hd__a21o_1 _07741_ (.A1(_02258_),
    .A2(_02260_),
    .B1(_02285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02293_));
 sky130_fd_sc_hd__clkbuf_1 _07742_ (.A(_02244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02294_));
 sky130_fd_sc_hd__and2_1 _07743_ (.A(_02199_),
    .B(_02252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02295_));
 sky130_fd_sc_hd__a21oi_1 _07744_ (.A1(_02181_),
    .A2(_02294_),
    .B1(_02295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02296_));
 sky130_fd_sc_hd__and3_1 _07745_ (.A(_02181_),
    .B(_02244_),
    .C(_02295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02297_));
 sky130_fd_sc_hd__nor2_1 _07746_ (.A(_02296_),
    .B(_02297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02298_));
 sky130_fd_sc_hd__nand2_1 _07747_ (.A(_02178_),
    .B(_02253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02299_));
 sky130_fd_sc_hd__xnor2_1 _07748_ (.A(_02298_),
    .B(_02299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02300_));
 sky130_fd_sc_hd__o21ba_1 _07749_ (.A1(_02275_),
    .A2(_02278_),
    .B1_N(_02276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02301_));
 sky130_fd_sc_hd__inv_2 _07750_ (.A(_02301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02302_));
 sky130_fd_sc_hd__xnor2_1 _07751_ (.A(_02300_),
    .B(_02302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02303_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07752_ (.A(_02253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02304_));
 sky130_fd_sc_hd__and2b_1 _07753_ (.A_N(_02280_),
    .B(_02279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02305_));
 sky130_fd_sc_hd__a31oi_1 _07754_ (.A1(_02165_),
    .A2(_02304_),
    .A3(_02281_),
    .B1(_02305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02306_));
 sky130_fd_sc_hd__nor2_1 _07755_ (.A(_02303_),
    .B(_02306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02307_));
 sky130_fd_sc_hd__and2_1 _07756_ (.A(_02303_),
    .B(_02306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02308_));
 sky130_fd_sc_hd__and2b_1 _07757_ (.A_N(_02282_),
    .B(_02283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02309_));
 sky130_fd_sc_hd__a21oi_1 _07758_ (.A1(_02255_),
    .A2(_02284_),
    .B1(_02309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02310_));
 sky130_fd_sc_hd__or3_1 _07759_ (.A(_02307_),
    .B(_02308_),
    .C(_02310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02311_));
 sky130_fd_sc_hd__nor2_1 _07760_ (.A(_02307_),
    .B(_02308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02312_));
 sky130_fd_sc_hd__or2b_1 _07761_ (.A(_02312_),
    .B_N(_02310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02313_));
 sky130_fd_sc_hd__nand2_1 _07762_ (.A(_02311_),
    .B(_02313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02314_));
 sky130_fd_sc_hd__a21oi_1 _07763_ (.A1(_02293_),
    .A2(_02289_),
    .B1(_02314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02315_));
 sky130_fd_sc_hd__and3_1 _07764_ (.A(_02293_),
    .B(_02289_),
    .C(_02314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02316_));
 sky130_fd_sc_hd__nor2_1 _07765_ (.A(_02315_),
    .B(_02316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02317_));
 sky130_fd_sc_hd__xor2_1 _07766_ (.A(_01813_),
    .B(_02317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02318_));
 sky130_fd_sc_hd__mux2_1 _07767_ (.A0(_02291_),
    .A1(_02318_),
    .S(_02240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02319_));
 sky130_fd_sc_hd__clkbuf_1 _07768_ (.A(_02319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[8] ));
 sky130_fd_sc_hd__a21o_1 _07769_ (.A1(_02293_),
    .A2(_02289_),
    .B1(_02314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02320_));
 sky130_fd_sc_hd__a31o_1 _07770_ (.A1(_02178_),
    .A2(_02304_),
    .A3(_02298_),
    .B1(_02297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02321_));
 sky130_fd_sc_hd__a22oi_1 _07771_ (.A1(_02252_),
    .A2(_02294_),
    .B1(_02304_),
    .B2(_02199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02322_));
 sky130_fd_sc_hd__and4_1 _07772_ (.A(_02199_),
    .B(_02252_),
    .C(_02294_),
    .D(_02253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02323_));
 sky130_fd_sc_hd__nor2_1 _07773_ (.A(_02322_),
    .B(_02323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02324_));
 sky130_fd_sc_hd__xnor2_1 _07774_ (.A(_02321_),
    .B(_02324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02325_));
 sky130_fd_sc_hd__a21oi_1 _07775_ (.A1(_02300_),
    .A2(_02302_),
    .B1(_02307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02326_));
 sky130_fd_sc_hd__xnor2_1 _07776_ (.A(_02325_),
    .B(_02326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02327_));
 sky130_fd_sc_hd__a21oi_1 _07777_ (.A1(_02311_),
    .A2(_02320_),
    .B1(_02327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02328_));
 sky130_fd_sc_hd__and3_1 _07778_ (.A(_02311_),
    .B(_02320_),
    .C(_02327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02329_));
 sky130_fd_sc_hd__or2_1 _07779_ (.A(_02328_),
    .B(_02329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02330_));
 sky130_fd_sc_hd__xnor2_1 _07780_ (.A(_01813_),
    .B(_02330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02331_));
 sky130_fd_sc_hd__mux2_1 _07781_ (.A0(_02318_),
    .A1(_02331_),
    .S(_02240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02332_));
 sky130_fd_sc_hd__clkbuf_1 _07782_ (.A(_02332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[9] ));
 sky130_fd_sc_hd__inv_2 _07783_ (.A(_02325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02333_));
 sky130_fd_sc_hd__a21o_1 _07784_ (.A1(_02307_),
    .A2(_02333_),
    .B1(_02328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02334_));
 sky130_fd_sc_hd__and3b_1 _07785_ (.A_N(_02295_),
    .B(_02304_),
    .C(_02294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02335_));
 sky130_fd_sc_hd__and2_1 _07786_ (.A(_02321_),
    .B(_02324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02336_));
 sky130_fd_sc_hd__and3_1 _07787_ (.A(_02300_),
    .B(_02302_),
    .C(_02333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02337_));
 sky130_fd_sc_hd__nor2_1 _07788_ (.A(_02336_),
    .B(_02337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02338_));
 sky130_fd_sc_hd__xnor2_1 _07789_ (.A(_02335_),
    .B(_02338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02339_));
 sky130_fd_sc_hd__xnor2_1 _07790_ (.A(_02334_),
    .B(_02339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02340_));
 sky130_fd_sc_hd__xnor2_1 _07791_ (.A(_01813_),
    .B(_02340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02341_));
 sky130_fd_sc_hd__mux2_1 _07792_ (.A0(_02331_),
    .A1(_02341_),
    .S(_02162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02342_));
 sky130_fd_sc_hd__clkbuf_1 _07793_ (.A(_02342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[10] ));
 sky130_fd_sc_hd__a22o_1 _07794_ (.A1(_02335_),
    .A2(_02337_),
    .B1(_02339_),
    .B2(_02334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02343_));
 sky130_fd_sc_hd__o211a_1 _07795_ (.A1(_02295_),
    .A2(_02336_),
    .B1(_02294_),
    .C1(_02304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02344_));
 sky130_fd_sc_hd__xnor2_1 _07796_ (.A(_01812_),
    .B(_02344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02345_));
 sky130_fd_sc_hd__xnor2_1 _07797_ (.A(_02343_),
    .B(_02345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02346_));
 sky130_fd_sc_hd__mux2_1 _07798_ (.A0(_02341_),
    .A1(_02346_),
    .S(_02162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02347_));
 sky130_fd_sc_hd__clkbuf_1 _07799_ (.A(_02347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[11] ));
 sky130_fd_sc_hd__mux2_1 _07800_ (.A0(_02346_),
    .A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._01_ ),
    .S(_02162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02348_));
 sky130_fd_sc_hd__clkbuf_1 _07801_ (.A(_02348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[12] ));
 sky130_fd_sc_hd__nand2_1 _07802_ (.A(_01275_),
    .B(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02349_));
 sky130_fd_sc_hd__xnor2_1 _07803_ (.A(_01274_),
    .B(_02349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[0] ));
 sky130_fd_sc_hd__and3_1 _07804_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[1] ),
    .B(_01288_),
    .C(_01290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02350_));
 sky130_fd_sc_hd__a21o_1 _07805_ (.A1(_01288_),
    .A2(_01290_),
    .B1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02351_));
 sky130_fd_sc_hd__or2b_1 _07806_ (.A(_02350_),
    .B_N(_02351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02352_));
 sky130_fd_sc_hd__nand2_1 _07807_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[0] ),
    .B(_01274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02353_));
 sky130_fd_sc_hd__xor2_1 _07808_ (.A(_02352_),
    .B(_02353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02354_));
 sky130_fd_sc_hd__mux2_1 _07809_ (.A0(_01291_),
    .A1(_02354_),
    .S(_01393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02355_));
 sky130_fd_sc_hd__clkbuf_1 _07810_ (.A(_02355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[1] ));
 sky130_fd_sc_hd__buf_2 _07811_ (.A(_01297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02356_));
 sky130_fd_sc_hd__a31o_1 _07812_ (.A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[0] ),
    .A2(_01274_),
    .A3(_02351_),
    .B1(_02350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02357_));
 sky130_fd_sc_hd__or2_1 _07813_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[2] ),
    .B(_01311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02358_));
 sky130_fd_sc_hd__nand2_1 _07814_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[2] ),
    .B(_01313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02359_));
 sky130_fd_sc_hd__nand3_1 _07815_ (.A(_02357_),
    .B(_02358_),
    .C(_02359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02360_));
 sky130_fd_sc_hd__a21o_1 _07816_ (.A1(_02358_),
    .A2(_02359_),
    .B1(_02357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02361_));
 sky130_fd_sc_hd__a31o_1 _07817_ (.A1(_02356_),
    .A2(_02360_),
    .A3(_02361_),
    .B1(_01319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[2] ));
 sky130_fd_sc_hd__nor2_1 _07818_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[3] ),
    .B(_01327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02362_));
 sky130_fd_sc_hd__and2_1 _07819_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[3] ),
    .B(_01327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02363_));
 sky130_fd_sc_hd__or2_1 _07820_ (.A(_02362_),
    .B(_02363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02364_));
 sky130_fd_sc_hd__and2_1 _07821_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[2] ),
    .B(_01313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02365_));
 sky130_fd_sc_hd__a21o_1 _07822_ (.A1(_02357_),
    .A2(_02358_),
    .B1(_02365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02366_));
 sky130_fd_sc_hd__xnor2_1 _07823_ (.A(_02364_),
    .B(_02366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02367_));
 sky130_fd_sc_hd__mux2_1 _07824_ (.A0(_01327_),
    .A1(_02367_),
    .S(_01393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02368_));
 sky130_fd_sc_hd__clkbuf_1 _07825_ (.A(_02368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[3] ));
 sky130_fd_sc_hd__xnor2_1 _07826_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[4] ),
    .B(_01341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02369_));
 sky130_fd_sc_hd__a221o_1 _07827_ (.A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[3] ),
    .A2(_01327_),
    .B1(_02357_),
    .B2(_02358_),
    .C1(_02365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02370_));
 sky130_fd_sc_hd__and2b_1 _07828_ (.A_N(_02362_),
    .B(_02370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02371_));
 sky130_fd_sc_hd__xnor2_1 _07829_ (.A(_02369_),
    .B(_02371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02372_));
 sky130_fd_sc_hd__mux2_1 _07830_ (.A0(_01341_),
    .A1(_02372_),
    .S(_01393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02373_));
 sky130_fd_sc_hd__clkbuf_1 _07831_ (.A(_02373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[4] ));
 sky130_fd_sc_hd__nand2_2 _07832_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[4] ),
    .B(_01341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02374_));
 sky130_fd_sc_hd__or3b_2 _07833_ (.A(_02362_),
    .B(_02369_),
    .C_N(_02370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02375_));
 sky130_fd_sc_hd__xnor2_2 _07834_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[5] ),
    .B(_01354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02376_));
 sky130_fd_sc_hd__nand3_1 _07835_ (.A(_02374_),
    .B(_02375_),
    .C(_02376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02377_));
 sky130_fd_sc_hd__a21o_1 _07836_ (.A1(_02374_),
    .A2(_02375_),
    .B1(_02376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02378_));
 sky130_fd_sc_hd__a31o_1 _07837_ (.A1(_02356_),
    .A2(_02377_),
    .A3(_02378_),
    .B1(_01364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[5] ));
 sky130_fd_sc_hd__xnor2_4 _07838_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[6] ),
    .B(_01367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02379_));
 sky130_fd_sc_hd__nand2_1 _07839_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[5] ),
    .B(_01354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02380_));
 sky130_fd_sc_hd__nor2_1 _07840_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[5] ),
    .B(_01354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02381_));
 sky130_fd_sc_hd__a31o_1 _07841_ (.A1(_02374_),
    .A2(_02375_),
    .A3(_02380_),
    .B1(_02381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02382_));
 sky130_fd_sc_hd__xor2_1 _07842_ (.A(_02379_),
    .B(_02382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02383_));
 sky130_fd_sc_hd__mux2_1 _07843_ (.A0(_01368_),
    .A1(_02383_),
    .S(_01393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02384_));
 sky130_fd_sc_hd__clkbuf_1 _07844_ (.A(_02384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[6] ));
 sky130_fd_sc_hd__a21oi_1 _07845_ (.A1(_01383_),
    .A2(_01384_),
    .B1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02385_));
 sky130_fd_sc_hd__and3_1 _07846_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[7] ),
    .B(_01383_),
    .C(_01384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02386_));
 sky130_fd_sc_hd__or2_2 _07847_ (.A(_02385_),
    .B(_02386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02387_));
 sky130_fd_sc_hd__nand2_1 _07848_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[6] ),
    .B(_01368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02388_));
 sky130_fd_sc_hd__o21ai_1 _07849_ (.A1(_02379_),
    .A2(_02382_),
    .B1(_02388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02389_));
 sky130_fd_sc_hd__xnor2_1 _07850_ (.A(_02387_),
    .B(_02389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02390_));
 sky130_fd_sc_hd__mux2_1 _07851_ (.A0(_01385_),
    .A1(_02390_),
    .S(_01392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02391_));
 sky130_fd_sc_hd__clkbuf_1 _07852_ (.A(_02391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[7] ));
 sky130_fd_sc_hd__and3_1 _07853_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[8] ),
    .B(_01398_),
    .C(_01399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02392_));
 sky130_fd_sc_hd__a21oi_1 _07854_ (.A1(_01398_),
    .A2(_01399_),
    .B1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02393_));
 sky130_fd_sc_hd__or2_1 _07855_ (.A(_02392_),
    .B(_02393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02394_));
 sky130_fd_sc_hd__and3b_1 _07856_ (.A_N(_02385_),
    .B(_01368_),
    .C(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02395_));
 sky130_fd_sc_hd__a2111oi_4 _07857_ (.A1(_02374_),
    .A2(_02380_),
    .B1(_02381_),
    .C1(_02379_),
    .D1(_02387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02396_));
 sky130_fd_sc_hd__nor4_2 _07858_ (.A(_02375_),
    .B(_02376_),
    .C(_02379_),
    .D(_02387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02397_));
 sky130_fd_sc_hd__nor4_2 _07859_ (.A(_02386_),
    .B(_02395_),
    .C(_02396_),
    .D(_02397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02398_));
 sky130_fd_sc_hd__xor2_1 _07860_ (.A(_02394_),
    .B(_02398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02399_));
 sky130_fd_sc_hd__mux2_1 _07861_ (.A0(_01401_),
    .A1(_02399_),
    .S(_01392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02400_));
 sky130_fd_sc_hd__clkbuf_1 _07862_ (.A(_02400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[8] ));
 sky130_fd_sc_hd__and3_1 _07863_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[9] ),
    .B(_01414_),
    .C(_01415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02401_));
 sky130_fd_sc_hd__a21oi_1 _07864_ (.A1(_01422_),
    .A2(_01415_),
    .B1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02402_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07865_ (.A(_02402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02403_));
 sky130_fd_sc_hd__o21ba_1 _07866_ (.A1(_02394_),
    .A2(_02398_),
    .B1_N(_02392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02404_));
 sky130_fd_sc_hd__o21ai_1 _07867_ (.A1(_02401_),
    .A2(_02403_),
    .B1(_02404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02405_));
 sky130_fd_sc_hd__o31a_1 _07868_ (.A1(_02401_),
    .A2(_02403_),
    .A3(_02404_),
    .B1(_01493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02406_));
 sky130_fd_sc_hd__a22o_1 _07869_ (.A1(_01371_),
    .A2(_01423_),
    .B1(_02405_),
    .B2(_02406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[9] ));
 sky130_fd_sc_hd__xnor2_2 _07870_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[10] ),
    .B(_01433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02407_));
 sky130_fd_sc_hd__nor2_1 _07871_ (.A(_02392_),
    .B(_02401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02408_));
 sky130_fd_sc_hd__o21a_1 _07872_ (.A1(_02394_),
    .A2(_02398_),
    .B1(_02408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02409_));
 sky130_fd_sc_hd__or3_1 _07873_ (.A(_02403_),
    .B(_02407_),
    .C(_02409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02410_));
 sky130_fd_sc_hd__o21ai_1 _07874_ (.A1(_02403_),
    .A2(_02409_),
    .B1(_02407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02411_));
 sky130_fd_sc_hd__a31o_1 _07875_ (.A1(_02356_),
    .A2(_02410_),
    .A3(_02411_),
    .B1(_01434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[10] ));
 sky130_fd_sc_hd__nand2_1 _07876_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[10] ),
    .B(_01433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02412_));
 sky130_fd_sc_hd__a21oi_1 _07877_ (.A1(_01439_),
    .A2(_01440_),
    .B1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02413_));
 sky130_fd_sc_hd__and3_1 _07878_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[11] ),
    .B(_01439_),
    .C(_01440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02414_));
 sky130_fd_sc_hd__or2_1 _07879_ (.A(_02413_),
    .B(_02414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02415_));
 sky130_fd_sc_hd__a21o_1 _07880_ (.A1(_02412_),
    .A2(_02410_),
    .B1(_02415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02416_));
 sky130_fd_sc_hd__nand3_1 _07881_ (.A(_02412_),
    .B(_02410_),
    .C(_02415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02417_));
 sky130_fd_sc_hd__a31o_1 _07882_ (.A1(_02356_),
    .A2(_02416_),
    .A3(_02417_),
    .B1(_01446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[11] ));
 sky130_fd_sc_hd__o21ba_1 _07883_ (.A1(_02412_),
    .A2(_02413_),
    .B1_N(_02414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02418_));
 sky130_fd_sc_hd__or4_1 _07884_ (.A(_02402_),
    .B(_02407_),
    .C(_02408_),
    .D(_02415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02419_));
 sky130_fd_sc_hd__or4_1 _07885_ (.A(_02392_),
    .B(_02393_),
    .C(_02401_),
    .D(_02402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02420_));
 sky130_fd_sc_hd__nor4_1 _07886_ (.A(_02407_),
    .B(_02420_),
    .C(_02413_),
    .D(_02414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02421_));
 sky130_fd_sc_hd__o41ai_2 _07887_ (.A1(_02386_),
    .A2(_02395_),
    .A3(_02396_),
    .A4(_02397_),
    .B1(_02421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02422_));
 sky130_fd_sc_hd__nand2_1 _07888_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[12] ),
    .B(_01455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02423_));
 sky130_fd_sc_hd__or2_1 _07889_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[12] ),
    .B(_01455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02424_));
 sky130_fd_sc_hd__nand2_1 _07890_ (.A(_02423_),
    .B(_02424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02425_));
 sky130_fd_sc_hd__a31o_1 _07891_ (.A1(_02418_),
    .A2(_02419_),
    .A3(_02422_),
    .B1(_02425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02426_));
 sky130_fd_sc_hd__or4_1 _07892_ (.A(_02403_),
    .B(_02407_),
    .C(_02409_),
    .D(_02415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02427_));
 sky130_fd_sc_hd__nand3_1 _07893_ (.A(_02425_),
    .B(_02418_),
    .C(_02427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02428_));
 sky130_fd_sc_hd__a31o_1 _07894_ (.A1(_02356_),
    .A2(_02426_),
    .A3(_02428_),
    .B1(_01462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[12] ));
 sky130_fd_sc_hd__and3_1 _07895_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[13] ),
    .B(_01463_),
    .C(_01466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02429_));
 sky130_fd_sc_hd__a21oi_1 _07896_ (.A1(_01463_),
    .A2(_01466_),
    .B1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02430_));
 sky130_fd_sc_hd__nor2_1 _07897_ (.A(_02429_),
    .B(_02430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02431_));
 sky130_fd_sc_hd__and2_1 _07898_ (.A(_02423_),
    .B(_02426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02432_));
 sky130_fd_sc_hd__xnor2_1 _07899_ (.A(_02431_),
    .B(_02432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02433_));
 sky130_fd_sc_hd__a21o_1 _07900_ (.A1(_01585_),
    .A2(_02433_),
    .B1(_01472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[13] ));
 sky130_fd_sc_hd__nand2_1 _07901_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[14] ),
    .B(_01476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02434_));
 sky130_fd_sc_hd__or2_1 _07902_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[14] ),
    .B(_01476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02435_));
 sky130_fd_sc_hd__nand2_1 _07903_ (.A(_02434_),
    .B(_02435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02436_));
 sky130_fd_sc_hd__nor2_1 _07904_ (.A(_02430_),
    .B(_02432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02437_));
 sky130_fd_sc_hd__nor2_1 _07905_ (.A(_02429_),
    .B(_02437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02438_));
 sky130_fd_sc_hd__or2_1 _07906_ (.A(_02436_),
    .B(_02438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02439_));
 sky130_fd_sc_hd__a21oi_1 _07907_ (.A1(_02436_),
    .A2(_02438_),
    .B1(_01371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02440_));
 sky130_fd_sc_hd__a21o_1 _07908_ (.A1(_02439_),
    .A2(_02440_),
    .B1(_01481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[14] ));
 sky130_fd_sc_hd__clkbuf_2 _07909_ (.A(_01297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02441_));
 sky130_fd_sc_hd__and2_1 _07910_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[15] ),
    .B(_01485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02442_));
 sky130_fd_sc_hd__nor2_1 _07911_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[15] ),
    .B(_01486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02443_));
 sky130_fd_sc_hd__or2_1 _07912_ (.A(_02442_),
    .B(_02443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02444_));
 sky130_fd_sc_hd__a21o_1 _07913_ (.A1(_02434_),
    .A2(_02439_),
    .B1(_02444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02445_));
 sky130_fd_sc_hd__nand3_1 _07914_ (.A(_02434_),
    .B(_02439_),
    .C(_02444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02446_));
 sky130_fd_sc_hd__a31o_1 _07915_ (.A1(_02441_),
    .A2(_02445_),
    .A3(_02446_),
    .B1(_01492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[15] ));
 sky130_fd_sc_hd__nor2_1 _07916_ (.A(_02436_),
    .B(_02444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02447_));
 sky130_fd_sc_hd__nand2_1 _07917_ (.A(_02431_),
    .B(_02447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02448_));
 sky130_fd_sc_hd__o21bai_1 _07918_ (.A1(_02423_),
    .A2(_02430_),
    .B1_N(_02429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02449_));
 sky130_fd_sc_hd__a22oi_1 _07919_ (.A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[15] ),
    .A2(_01486_),
    .B1(_02447_),
    .B2(_02449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02450_));
 sky130_fd_sc_hd__o221a_2 _07920_ (.A1(_02434_),
    .A2(_02443_),
    .B1(_02448_),
    .B2(_02426_),
    .C1(_02450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02451_));
 sky130_fd_sc_hd__nand2_1 _07921_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[16] ),
    .B(_01503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02452_));
 sky130_fd_sc_hd__or2_1 _07922_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[16] ),
    .B(_01505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02453_));
 sky130_fd_sc_hd__nand2_1 _07923_ (.A(_02452_),
    .B(_02453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02454_));
 sky130_fd_sc_hd__or2_1 _07924_ (.A(_02451_),
    .B(_02454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02455_));
 sky130_fd_sc_hd__nand2_1 _07925_ (.A(_02451_),
    .B(_02454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02456_));
 sky130_fd_sc_hd__a31o_1 _07926_ (.A1(_02441_),
    .A2(_02455_),
    .A3(_02456_),
    .B1(_01584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[16] ));
 sky130_fd_sc_hd__o21a_1 _07927_ (.A1(_02451_),
    .A2(_02454_),
    .B1(_02452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02457_));
 sky130_fd_sc_hd__nand2_1 _07928_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[17] ),
    .B(_01521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02458_));
 sky130_fd_sc_hd__or2_1 _07929_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[17] ),
    .B(_01502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02459_));
 sky130_fd_sc_hd__nand2_1 _07930_ (.A(_02458_),
    .B(_02459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02460_));
 sky130_fd_sc_hd__xor2_1 _07931_ (.A(_02457_),
    .B(_02460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02461_));
 sky130_fd_sc_hd__clkbuf_2 _07932_ (.A(_01516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02462_));
 sky130_fd_sc_hd__a21o_1 _07933_ (.A1(_01585_),
    .A2(_02461_),
    .B1(_02462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[17] ));
 sky130_fd_sc_hd__or2b_1 _07934_ (.A(_02457_),
    .B_N(_02459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02463_));
 sky130_fd_sc_hd__nand2_1 _07935_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[18] ),
    .B(_01503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02464_));
 sky130_fd_sc_hd__or2_1 _07936_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[18] ),
    .B(_01505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02465_));
 sky130_fd_sc_hd__nand2_1 _07937_ (.A(_02464_),
    .B(_02465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02466_));
 sky130_fd_sc_hd__a21o_1 _07938_ (.A1(_02458_),
    .A2(_02463_),
    .B1(_02466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02467_));
 sky130_fd_sc_hd__nand3_1 _07939_ (.A(_02458_),
    .B(_02463_),
    .C(_02466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02468_));
 sky130_fd_sc_hd__clkbuf_2 _07940_ (.A(_01515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02469_));
 sky130_fd_sc_hd__a31o_1 _07941_ (.A1(_02441_),
    .A2(_02467_),
    .A3(_02468_),
    .B1(_02469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[18] ));
 sky130_fd_sc_hd__xnor2_1 _07942_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[19] ),
    .B(_01509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02470_));
 sky130_fd_sc_hd__a21o_1 _07943_ (.A1(_02464_),
    .A2(_02467_),
    .B1(_02470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02471_));
 sky130_fd_sc_hd__nand3_1 _07944_ (.A(_02464_),
    .B(_02467_),
    .C(_02470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02472_));
 sky130_fd_sc_hd__a31o_1 _07945_ (.A1(_02441_),
    .A2(_02471_),
    .A3(_02472_),
    .B1(_02469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[19] ));
 sky130_fd_sc_hd__nand2_1 _07946_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[20] ),
    .B(_01503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02473_));
 sky130_fd_sc_hd__or2_1 _07947_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[20] ),
    .B(_01505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02474_));
 sky130_fd_sc_hd__nand2_1 _07948_ (.A(_02473_),
    .B(_02474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02475_));
 sky130_fd_sc_hd__or4_1 _07949_ (.A(_02454_),
    .B(_02460_),
    .C(_02466_),
    .D(_02470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02476_));
 sky130_fd_sc_hd__o41a_1 _07950_ (.A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[16] ),
    .A2(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[17] ),
    .A3(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[18] ),
    .A4(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[19] ),
    .B1(_01511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02477_));
 sky130_fd_sc_hd__o21ba_1 _07951_ (.A1(_02451_),
    .A2(_02476_),
    .B1_N(_02477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02478_));
 sky130_fd_sc_hd__or2_1 _07952_ (.A(_02475_),
    .B(_02478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02479_));
 sky130_fd_sc_hd__nand2_1 _07953_ (.A(_02475_),
    .B(_02478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02480_));
 sky130_fd_sc_hd__a31o_1 _07954_ (.A1(_02441_),
    .A2(_02479_),
    .A3(_02480_),
    .B1(_02469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[20] ));
 sky130_fd_sc_hd__nand2_1 _07955_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[21] ),
    .B(_01503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02481_));
 sky130_fd_sc_hd__or2_1 _07956_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[21] ),
    .B(_01521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02482_));
 sky130_fd_sc_hd__nand2_1 _07957_ (.A(_02481_),
    .B(_02482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02483_));
 sky130_fd_sc_hd__a21o_1 _07958_ (.A1(_02473_),
    .A2(_02479_),
    .B1(_02483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02484_));
 sky130_fd_sc_hd__a31oi_1 _07959_ (.A1(_02473_),
    .A2(_02479_),
    .A3(_02483_),
    .B1(_01371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02485_));
 sky130_fd_sc_hd__a21o_1 _07960_ (.A1(_02484_),
    .A2(_02485_),
    .B1(_02462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[21] ));
 sky130_fd_sc_hd__a21bo_1 _07961_ (.A1(_02473_),
    .A2(_02479_),
    .B1_N(_02482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02486_));
 sky130_fd_sc_hd__and2_1 _07962_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[22] ),
    .B(_01502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02487_));
 sky130_fd_sc_hd__nor2_1 _07963_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[22] ),
    .B(_01521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02488_));
 sky130_fd_sc_hd__or2_1 _07964_ (.A(_02487_),
    .B(_02488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02489_));
 sky130_fd_sc_hd__a21oi_1 _07965_ (.A1(_02481_),
    .A2(_02486_),
    .B1(_02489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02490_));
 sky130_fd_sc_hd__a31o_1 _07966_ (.A1(_02481_),
    .A2(_02486_),
    .A3(_02489_),
    .B1(_01460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02491_));
 sky130_fd_sc_hd__o21bai_1 _07967_ (.A1(_02490_),
    .A2(_02491_),
    .B1_N(_01546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[22] ));
 sky130_fd_sc_hd__xor2_1 _07968_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[23] ),
    .B(_01509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02492_));
 sky130_fd_sc_hd__o21ai_1 _07969_ (.A1(_02487_),
    .A2(_02490_),
    .B1(_02492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02493_));
 sky130_fd_sc_hd__or3_1 _07970_ (.A(_02487_),
    .B(_02490_),
    .C(_02492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02494_));
 sky130_fd_sc_hd__a31o_1 _07971_ (.A1(_01407_),
    .A2(_02493_),
    .A3(_02494_),
    .B1(_02469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[23] ));
 sky130_fd_sc_hd__or4b_1 _07972_ (.A(_02475_),
    .B(_02483_),
    .C(_02489_),
    .D_N(_02492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02495_));
 sky130_fd_sc_hd__or2_1 _07973_ (.A(_02476_),
    .B(_02495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02496_));
 sky130_fd_sc_hd__o41a_1 _07974_ (.A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[20] ),
    .A2(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[21] ),
    .A3(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[22] ),
    .A4(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[23] ),
    .B1(_01566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02497_));
 sky130_fd_sc_hd__nor2_1 _07975_ (.A(_02477_),
    .B(_02497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02498_));
 sky130_fd_sc_hd__o21ai_4 _07976_ (.A1(_02451_),
    .A2(_02496_),
    .B1(_02498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02499_));
 sky130_fd_sc_hd__xor2_1 _07977_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[24] ),
    .B(_01566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02500_));
 sky130_fd_sc_hd__nand2_1 _07978_ (.A(_02499_),
    .B(_02500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02501_));
 sky130_fd_sc_hd__o21a_1 _07979_ (.A1(_02499_),
    .A2(_02500_),
    .B1(_01493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02502_));
 sky130_fd_sc_hd__a21o_1 _07980_ (.A1(_02501_),
    .A2(_02502_),
    .B1(_02462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[24] ));
 sky130_fd_sc_hd__xor2_1 _07981_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[25] ),
    .B(_01566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02503_));
 sky130_fd_sc_hd__a22o_1 _07982_ (.A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[24] ),
    .A2(_01573_),
    .B1(_02499_),
    .B2(_02500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02504_));
 sky130_fd_sc_hd__xor2_1 _07983_ (.A(_02503_),
    .B(_02504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02505_));
 sky130_fd_sc_hd__a21o_1 _07984_ (.A1(_01585_),
    .A2(_02505_),
    .B1(_02462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[25] ));
 sky130_fd_sc_hd__o21ai_1 _07985_ (.A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[24] ),
    .A2(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[25] ),
    .B1(_01514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02506_));
 sky130_fd_sc_hd__and2_1 _07986_ (.A(_02500_),
    .B(_02503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02507_));
 sky130_fd_sc_hd__nand2_1 _07987_ (.A(_02499_),
    .B(_02507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02508_));
 sky130_fd_sc_hd__nand2_1 _07988_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[26] ),
    .B(_01541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02509_));
 sky130_fd_sc_hd__or2_1 _07989_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[26] ),
    .B(_01511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02510_));
 sky130_fd_sc_hd__nand2_1 _07990_ (.A(_02509_),
    .B(_02510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02511_));
 sky130_fd_sc_hd__a21o_1 _07991_ (.A1(_02506_),
    .A2(_02508_),
    .B1(_02511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02512_));
 sky130_fd_sc_hd__nand3_1 _07992_ (.A(_02511_),
    .B(_02506_),
    .C(_02508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02513_));
 sky130_fd_sc_hd__a31o_1 _07993_ (.A1(_01407_),
    .A2(_02512_),
    .A3(_02513_),
    .B1(_02469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[26] ));
 sky130_fd_sc_hd__xnor2_1 _07994_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[27] ),
    .B(_01512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02514_));
 sky130_fd_sc_hd__nand2_1 _07995_ (.A(_02509_),
    .B(_02512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02515_));
 sky130_fd_sc_hd__xnor2_1 _07996_ (.A(_02514_),
    .B(_02515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02516_));
 sky130_fd_sc_hd__a21o_1 _07997_ (.A1(_01585_),
    .A2(_02516_),
    .B1(_02462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[27] ));
 sky130_fd_sc_hd__nor2_1 _07998_ (.A(_02511_),
    .B(_02514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02517_));
 sky130_fd_sc_hd__o41a_1 _07999_ (.A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[24] ),
    .A2(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[25] ),
    .A3(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[26] ),
    .A4(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[27] ),
    .B1(_01571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02518_));
 sky130_fd_sc_hd__a31oi_2 _08000_ (.A1(_02499_),
    .A2(_02507_),
    .A3(_02517_),
    .B1(_02518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02519_));
 sky130_fd_sc_hd__and2_1 _08001_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[28] ),
    .B(_01512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02520_));
 sky130_fd_sc_hd__nor2_1 _08002_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[28] ),
    .B(_01571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02521_));
 sky130_fd_sc_hd__or2_1 _08003_ (.A(_02520_),
    .B(_02521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02522_));
 sky130_fd_sc_hd__nor2_1 _08004_ (.A(_02519_),
    .B(_02522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02523_));
 sky130_fd_sc_hd__a21o_1 _08005_ (.A1(_02519_),
    .A2(_02522_),
    .B1(_01460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02524_));
 sky130_fd_sc_hd__o21bai_1 _08006_ (.A1(_02523_),
    .A2(_02524_),
    .B1_N(_01516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[28] ));
 sky130_fd_sc_hd__nand2_1 _08007_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[29] ),
    .B(_01513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02525_));
 sky130_fd_sc_hd__or2_1 _08008_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[29] ),
    .B(_01513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02526_));
 sky130_fd_sc_hd__o211ai_1 _08009_ (.A1(_02520_),
    .A2(_02523_),
    .B1(_02525_),
    .C1(_02526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02527_));
 sky130_fd_sc_hd__a211o_1 _08010_ (.A1(_02525_),
    .A2(_02526_),
    .B1(_02520_),
    .C1(_02523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02528_));
 sky130_fd_sc_hd__a31o_1 _08011_ (.A1(_01407_),
    .A2(_02527_),
    .A3(_02528_),
    .B1(_01546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[29] ));
 sky130_fd_sc_hd__o21ai_1 _08012_ (.A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[28] ),
    .A2(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[29] ),
    .B1(_01514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02529_));
 sky130_fd_sc_hd__or4bb_1 _08013_ (.A(_02519_),
    .B(_02522_),
    .C_N(_02525_),
    .D_N(_02526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02530_));
 sky130_fd_sc_hd__nand2_1 _08014_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[30] ),
    .B(_01572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02531_));
 sky130_fd_sc_hd__or2_1 _08015_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[30] ),
    .B(_01572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02532_));
 sky130_fd_sc_hd__nand2_1 _08016_ (.A(_02531_),
    .B(_02532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02533_));
 sky130_fd_sc_hd__a21o_1 _08017_ (.A1(_02529_),
    .A2(_02530_),
    .B1(_02533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02534_));
 sky130_fd_sc_hd__nand3_1 _08018_ (.A(_02533_),
    .B(_02529_),
    .C(_02530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02535_));
 sky130_fd_sc_hd__a31o_1 _08019_ (.A1(_01407_),
    .A2(_02534_),
    .A3(_02535_),
    .B1(_01546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[30] ));
 sky130_fd_sc_hd__xnor2_1 _08020_ (.A(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[31] ),
    .B(_01573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02536_));
 sky130_fd_sc_hd__a21oi_1 _08021_ (.A1(_02531_),
    .A2(_02534_),
    .B1(_02536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02537_));
 sky130_fd_sc_hd__a31o_1 _08022_ (.A1(_02531_),
    .A2(_02534_),
    .A3(_02536_),
    .B1(_01318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02538_));
 sky130_fd_sc_hd__o21bai_1 _08023_ (.A1(_02537_),
    .A2(_02538_),
    .B1_N(_01516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[31] ));
 sky130_fd_sc_hd__buf_2 _08024_ (.A(\sa_inst.sak._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02539_));
 sky130_fd_sc_hd__clkbuf_4 _08025_ (.A(_02539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02540_));
 sky130_fd_sc_hd__mux2_1 _08026_ (.A0(\sa_inst.sak._40_[0] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[0] ),
    .S(_02540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02541_));
 sky130_fd_sc_hd__clkbuf_1 _08027_ (.A(_02541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ));
 sky130_fd_sc_hd__mux2_1 _08028_ (.A0(\sa_inst.sak._40_[1] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[1] ),
    .S(_02540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02542_));
 sky130_fd_sc_hd__clkbuf_1 _08029_ (.A(_02542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ));
 sky130_fd_sc_hd__clkbuf_4 _08030_ (.A(\sa_inst.sak._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02543_));
 sky130_fd_sc_hd__clkbuf_2 _08031_ (.A(_02543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02544_));
 sky130_fd_sc_hd__mux2_1 _08032_ (.A0(\sa_inst.sak._40_[2] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[2] ),
    .S(_02544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02545_));
 sky130_fd_sc_hd__clkbuf_1 _08033_ (.A(_02545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ));
 sky130_fd_sc_hd__mux2_1 _08034_ (.A0(\sa_inst.sak._40_[3] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[3] ),
    .S(_02544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02546_));
 sky130_fd_sc_hd__clkbuf_1 _08035_ (.A(_02546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ));
 sky130_fd_sc_hd__mux2_1 _08036_ (.A0(\sa_inst.sak._40_[4] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[4] ),
    .S(_02544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02547_));
 sky130_fd_sc_hd__clkbuf_1 _08037_ (.A(_02547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ));
 sky130_fd_sc_hd__mux2_1 _08038_ (.A0(\sa_inst.sak._40_[5] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[5] ),
    .S(_02544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02548_));
 sky130_fd_sc_hd__clkbuf_1 _08039_ (.A(_02548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ));
 sky130_fd_sc_hd__mux2_1 _08040_ (.A0(\sa_inst.sak._40_[6] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[6] ),
    .S(_02544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02549_));
 sky130_fd_sc_hd__clkbuf_1 _08041_ (.A(_02549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ));
 sky130_fd_sc_hd__clkbuf_2 _08042_ (.A(_02543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02550_));
 sky130_fd_sc_hd__mux2_1 _08043_ (.A0(\sa_inst.sak._40_[7] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[7] ),
    .S(_02550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02551_));
 sky130_fd_sc_hd__clkbuf_1 _08044_ (.A(_02551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ));
 sky130_fd_sc_hd__mux2_1 _08045_ (.A0(\sa_inst.sak._40_[8] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[8] ),
    .S(_02550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02552_));
 sky130_fd_sc_hd__clkbuf_1 _08046_ (.A(_02552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ));
 sky130_fd_sc_hd__mux2_1 _08047_ (.A0(\sa_inst.sak._40_[9] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[9] ),
    .S(_02550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02553_));
 sky130_fd_sc_hd__clkbuf_1 _08048_ (.A(_02553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ));
 sky130_fd_sc_hd__mux2_1 _08049_ (.A0(\sa_inst.sak._40_[10] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[10] ),
    .S(_02550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02554_));
 sky130_fd_sc_hd__clkbuf_1 _08050_ (.A(_02554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ));
 sky130_fd_sc_hd__mux2_1 _08051_ (.A0(\sa_inst.sak._40_[11] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[11] ),
    .S(_02550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02555_));
 sky130_fd_sc_hd__clkbuf_1 _08052_ (.A(_02555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ));
 sky130_fd_sc_hd__buf_2 _08053_ (.A(_02543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02556_));
 sky130_fd_sc_hd__mux2_1 _08054_ (.A0(\sa_inst.sak._40_[12] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[12] ),
    .S(_02556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02557_));
 sky130_fd_sc_hd__clkbuf_1 _08055_ (.A(_02557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ));
 sky130_fd_sc_hd__mux2_1 _08056_ (.A0(\sa_inst.sak._40_[13] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[13] ),
    .S(_02556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02558_));
 sky130_fd_sc_hd__clkbuf_1 _08057_ (.A(_02558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ));
 sky130_fd_sc_hd__mux2_1 _08058_ (.A0(\sa_inst.sak._40_[14] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[14] ),
    .S(_02556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02559_));
 sky130_fd_sc_hd__clkbuf_1 _08059_ (.A(_02559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ));
 sky130_fd_sc_hd__mux2_1 _08060_ (.A0(\sa_inst.sak._40_[15] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[15] ),
    .S(_02556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02560_));
 sky130_fd_sc_hd__clkbuf_1 _08061_ (.A(_02560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ));
 sky130_fd_sc_hd__mux2_1 _08062_ (.A0(\sa_inst.sak._40_[16] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[16] ),
    .S(_02556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02561_));
 sky130_fd_sc_hd__clkbuf_1 _08063_ (.A(_02561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ));
 sky130_fd_sc_hd__clkbuf_2 _08064_ (.A(_02539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02562_));
 sky130_fd_sc_hd__mux2_1 _08065_ (.A0(\sa_inst.sak._40_[17] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[17] ),
    .S(_02562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02563_));
 sky130_fd_sc_hd__clkbuf_1 _08066_ (.A(_02563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ));
 sky130_fd_sc_hd__mux2_1 _08067_ (.A0(\sa_inst.sak._40_[18] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[18] ),
    .S(_02562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02564_));
 sky130_fd_sc_hd__clkbuf_1 _08068_ (.A(_02564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ));
 sky130_fd_sc_hd__mux2_1 _08069_ (.A0(\sa_inst.sak._40_[19] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[19] ),
    .S(_02562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02565_));
 sky130_fd_sc_hd__clkbuf_1 _08070_ (.A(_02565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ));
 sky130_fd_sc_hd__mux2_1 _08071_ (.A0(\sa_inst.sak._40_[20] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[20] ),
    .S(_02562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02566_));
 sky130_fd_sc_hd__clkbuf_1 _08072_ (.A(_02566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ));
 sky130_fd_sc_hd__mux2_1 _08073_ (.A0(\sa_inst.sak._40_[21] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[21] ),
    .S(_02562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02567_));
 sky130_fd_sc_hd__clkbuf_1 _08074_ (.A(_02567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ));
 sky130_fd_sc_hd__buf_2 _08075_ (.A(_02539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02568_));
 sky130_fd_sc_hd__mux2_1 _08076_ (.A0(\sa_inst.sak._40_[22] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[22] ),
    .S(_02568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02569_));
 sky130_fd_sc_hd__clkbuf_1 _08077_ (.A(_02569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ));
 sky130_fd_sc_hd__mux2_1 _08078_ (.A0(\sa_inst.sak._40_[23] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[23] ),
    .S(_02568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02570_));
 sky130_fd_sc_hd__clkbuf_1 _08079_ (.A(_02570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ));
 sky130_fd_sc_hd__mux2_1 _08080_ (.A0(\sa_inst.sak._40_[24] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[24] ),
    .S(_02568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02571_));
 sky130_fd_sc_hd__clkbuf_1 _08081_ (.A(_02571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ));
 sky130_fd_sc_hd__mux2_1 _08082_ (.A0(\sa_inst.sak._40_[25] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[25] ),
    .S(_02568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02572_));
 sky130_fd_sc_hd__clkbuf_1 _08083_ (.A(_02572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ));
 sky130_fd_sc_hd__mux2_1 _08084_ (.A0(\sa_inst.sak._40_[26] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[26] ),
    .S(_02568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02573_));
 sky130_fd_sc_hd__clkbuf_1 _08085_ (.A(_02573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ));
 sky130_fd_sc_hd__buf_2 _08086_ (.A(_02539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02574_));
 sky130_fd_sc_hd__mux2_1 _08087_ (.A0(\sa_inst.sak._40_[27] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[27] ),
    .S(_02574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02575_));
 sky130_fd_sc_hd__clkbuf_1 _08088_ (.A(_02575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ));
 sky130_fd_sc_hd__mux2_1 _08089_ (.A0(\sa_inst.sak._40_[28] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[28] ),
    .S(_02574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02576_));
 sky130_fd_sc_hd__clkbuf_1 _08090_ (.A(_02576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ));
 sky130_fd_sc_hd__mux2_1 _08091_ (.A0(\sa_inst.sak._40_[29] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[29] ),
    .S(_02574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02577_));
 sky130_fd_sc_hd__clkbuf_1 _08092_ (.A(_02577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ));
 sky130_fd_sc_hd__mux2_1 _08093_ (.A0(\sa_inst.sak._40_[30] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[30] ),
    .S(_02574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02578_));
 sky130_fd_sc_hd__clkbuf_1 _08094_ (.A(_02578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ));
 sky130_fd_sc_hd__mux2_1 _08095_ (.A0(\sa_inst.sak._40_[31] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[31] ),
    .S(_02574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02579_));
 sky130_fd_sc_hd__clkbuf_1 _08096_ (.A(_02579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ));
 sky130_fd_sc_hd__clkbuf_2 _08097_ (.A(_02539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02580_));
 sky130_fd_sc_hd__mux2_1 _08098_ (.A0(\sa_inst.sak._40_[32] ),
    .A1(\sa_inst.sak.rows:2.cols:1.pe_ij._02_ ),
    .S(_02580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02581_));
 sky130_fd_sc_hd__clkbuf_1 _08099_ (.A(_02581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ));
 sky130_fd_sc_hd__inv_2 _08100_ (.A(\sa_inst.sak._13_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02582_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08101_ (.A(_02582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02583_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08102_ (.A(_02583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02584_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08103_ (.A(\sa_inst.sak._13_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02585_));
 sky130_fd_sc_hd__inv_2 _08104_ (.A(_02585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02586_));
 sky130_fd_sc_hd__clkbuf_2 _08105_ (.A(\sa_inst.sak._13_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02587_));
 sky130_fd_sc_hd__mux4_2 _08106_ (.A0(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .A2(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .A3(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .S0(\sa_inst.sak._13_[0] ),
    .S1(_02587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02588_));
 sky130_fd_sc_hd__clkbuf_2 _08107_ (.A(\sa_inst.sak._13_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02589_));
 sky130_fd_sc_hd__mux2_1 _08108_ (.A0(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ),
    .A1(\sa_inst.sak._13_[4] ),
    .S(_02589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02590_));
 sky130_fd_sc_hd__and2b_1 _08109_ (.A_N(_02587_),
    .B(_02585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02591_));
 sky130_fd_sc_hd__a22o_1 _08110_ (.A1(_02586_),
    .A2(_02588_),
    .B1(_02590_),
    .B2(_02591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02592_));
 sky130_fd_sc_hd__nand2_1 _08111_ (.A(_02584_),
    .B(_02592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02593_));
 sky130_fd_sc_hd__nand2_1 _08112_ (.A(_01828_),
    .B(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02594_));
 sky130_fd_sc_hd__xor2_1 _08113_ (.A(_02593_),
    .B(_02594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[0] ));
 sky130_fd_sc_hd__or2b_1 _08114_ (.A(_02587_),
    .B_N(\sa_inst.sak._13_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02595_));
 sky130_fd_sc_hd__clkbuf_2 _08115_ (.A(\sa_inst.sak._13_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02596_));
 sky130_fd_sc_hd__or2b_1 _08116_ (.A(_02596_),
    .B_N(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02597_));
 sky130_fd_sc_hd__mux4_2 _08117_ (.A0(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .A2(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .A3(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .S0(_02589_),
    .S1(_02587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02598_));
 sky130_fd_sc_hd__a2bb2o_1 _08118_ (.A1_N(_02595_),
    .A2_N(_02597_),
    .B1(_02598_),
    .B2(_02586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02599_));
 sky130_fd_sc_hd__and3_1 _08119_ (.A(_02582_),
    .B(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[0] ),
    .C(_02592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02600_));
 sky130_fd_sc_hd__and3_1 _08120_ (.A(_02582_),
    .B(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[1] ),
    .C(_02599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02601_));
 sky130_fd_sc_hd__a21o_1 _08121_ (.A1(_02583_),
    .A2(_02599_),
    .B1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02602_));
 sky130_fd_sc_hd__or2b_1 _08122_ (.A(_02601_),
    .B_N(_02602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02603_));
 sky130_fd_sc_hd__xnor2_1 _08123_ (.A(_02600_),
    .B(_02603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02604_));
 sky130_fd_sc_hd__and2_1 _08124_ (.A(_01826_),
    .B(_02604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02605_));
 sky130_fd_sc_hd__a31o_1 _08125_ (.A1(_01911_),
    .A2(_02584_),
    .A3(_02599_),
    .B1(_02605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[1] ));
 sky130_fd_sc_hd__mux2_1 _08126_ (.A0(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .S(\sa_inst.sak._13_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02606_));
 sky130_fd_sc_hd__and2_1 _08127_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .B(_02589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02607_));
 sky130_fd_sc_hd__and2b_1 _08128_ (.A_N(_02589_),
    .B(\sa_inst.sak._13_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02608_));
 sky130_fd_sc_hd__mux2_1 _08129_ (.A0(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ),
    .S(\sa_inst.sak._13_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02609_));
 sky130_fd_sc_hd__inv_2 _08130_ (.A(\sa_inst.sak._13_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02610_));
 sky130_fd_sc_hd__mux4_1 _08131_ (.A0(_02606_),
    .A1(_02607_),
    .A2(_02608_),
    .A3(_02609_),
    .S0(_02610_),
    .S1(_02585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02611_));
 sky130_fd_sc_hd__and2_1 _08132_ (.A(_02582_),
    .B(_02611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02612_));
 sky130_fd_sc_hd__a21o_1 _08133_ (.A1(_02600_),
    .A2(_02602_),
    .B1(_02601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02613_));
 sky130_fd_sc_hd__or2_1 _08134_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[2] ),
    .B(_02612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02614_));
 sky130_fd_sc_hd__nand2_1 _08135_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[2] ),
    .B(_02612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02615_));
 sky130_fd_sc_hd__nand2_1 _08136_ (.A(_02614_),
    .B(_02615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02616_));
 sky130_fd_sc_hd__xnor2_1 _08137_ (.A(_02613_),
    .B(_02616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02617_));
 sky130_fd_sc_hd__buf_2 _08138_ (.A(_01825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02618_));
 sky130_fd_sc_hd__mux2_1 _08139_ (.A0(_02612_),
    .A1(_02617_),
    .S(_02618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02619_));
 sky130_fd_sc_hd__clkbuf_1 _08140_ (.A(_02619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[2] ));
 sky130_fd_sc_hd__mux2_1 _08141_ (.A0(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .S(_02596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02620_));
 sky130_fd_sc_hd__clkbuf_2 _08142_ (.A(_02589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02621_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08143_ (.A(_02587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02622_));
 sky130_fd_sc_hd__a21o_1 _08144_ (.A1(_02621_),
    .A2(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .B1(_02622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02623_));
 sky130_fd_sc_hd__o211a_1 _08145_ (.A1(_02610_),
    .A2(_02620_),
    .B1(_02623_),
    .C1(_02586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02624_));
 sky130_fd_sc_hd__mux2_1 _08146_ (.A0(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ),
    .S(_02596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02625_));
 sky130_fd_sc_hd__and2_1 _08147_ (.A(_02591_),
    .B(_02625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02626_));
 sky130_fd_sc_hd__o21a_1 _08148_ (.A1(_02624_),
    .A2(_02626_),
    .B1(_02583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02627_));
 sky130_fd_sc_hd__nor2_1 _08149_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[3] ),
    .B(_02627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02628_));
 sky130_fd_sc_hd__and2_1 _08150_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[3] ),
    .B(_02627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02629_));
 sky130_fd_sc_hd__or2_1 _08151_ (.A(_02628_),
    .B(_02629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02630_));
 sky130_fd_sc_hd__and3_1 _08152_ (.A(_02584_),
    .B(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[2] ),
    .C(_02611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02631_));
 sky130_fd_sc_hd__a21o_1 _08153_ (.A1(_02613_),
    .A2(_02614_),
    .B1(_02631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02632_));
 sky130_fd_sc_hd__xnor2_1 _08154_ (.A(_02630_),
    .B(_02632_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02633_));
 sky130_fd_sc_hd__mux2_1 _08155_ (.A0(_02627_),
    .A1(_02633_),
    .S(_02618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02634_));
 sky130_fd_sc_hd__clkbuf_1 _08156_ (.A(_02634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[3] ));
 sky130_fd_sc_hd__buf_4 _08157_ (.A(_01850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02635_));
 sky130_fd_sc_hd__mux2_1 _08158_ (.A0(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .S(_02596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02636_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08159_ (.A(_02585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02637_));
 sky130_fd_sc_hd__a21o_1 _08160_ (.A1(_02622_),
    .A2(_02636_),
    .B1(_02637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02638_));
 sky130_fd_sc_hd__mux2_1 _08161_ (.A0(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .S(_02596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02639_));
 sky130_fd_sc_hd__nand2_1 _08162_ (.A(_02622_),
    .B(_02585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02640_));
 sky130_fd_sc_hd__o22a_1 _08163_ (.A1(_02639_),
    .A2(_02595_),
    .B1(_02640_),
    .B2(_02590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02641_));
 sky130_fd_sc_hd__and3_1 _08164_ (.A(_02582_),
    .B(_02638_),
    .C(_02641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02642_));
 sky130_fd_sc_hd__nand2_1 _08165_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[4] ),
    .B(_02642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02643_));
 sky130_fd_sc_hd__or2_1 _08166_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[4] ),
    .B(_02642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02644_));
 sky130_fd_sc_hd__nand2_1 _08167_ (.A(_02643_),
    .B(_02644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02645_));
 sky130_fd_sc_hd__a211oi_1 _08168_ (.A1(_02613_),
    .A2(_02614_),
    .B1(_02631_),
    .C1(_02629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02646_));
 sky130_fd_sc_hd__or2_1 _08169_ (.A(_02628_),
    .B(_02646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02647_));
 sky130_fd_sc_hd__or2_1 _08170_ (.A(_02645_),
    .B(_02647_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02648_));
 sky130_fd_sc_hd__a21oi_1 _08171_ (.A1(_02645_),
    .A2(_02647_),
    .B1(_01924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02649_));
 sky130_fd_sc_hd__a22o_1 _08172_ (.A1(_02635_),
    .A2(_02642_),
    .B1(_02648_),
    .B2(_02649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[4] ));
 sky130_fd_sc_hd__mux2_1 _08173_ (.A0(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .S(_02621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02650_));
 sky130_fd_sc_hd__mux2_1 _08174_ (.A0(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .S(_02621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02651_));
 sky130_fd_sc_hd__a21o_1 _08175_ (.A1(_02622_),
    .A2(_02651_),
    .B1(_02637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02652_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08176_ (.A(_02622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02653_));
 sky130_fd_sc_hd__clkbuf_2 _08177_ (.A(_02637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02654_));
 sky130_fd_sc_hd__a31oi_1 _08178_ (.A1(_02653_),
    .A2(_02654_),
    .A3(_02597_),
    .B1(\sa_inst.sak._13_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02655_));
 sky130_fd_sc_hd__o211a_2 _08179_ (.A1(_02595_),
    .A2(_02650_),
    .B1(_02652_),
    .C1(_02655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02656_));
 sky130_fd_sc_hd__xnor2_1 _08180_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[5] ),
    .B(_02656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02657_));
 sky130_fd_sc_hd__a31o_1 _08181_ (.A1(_02643_),
    .A2(_02648_),
    .A3(_02657_),
    .B1(_01910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02658_));
 sky130_fd_sc_hd__a21oi_1 _08182_ (.A1(_02643_),
    .A2(_02648_),
    .B1(_02657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02659_));
 sky130_fd_sc_hd__a2bb2o_1 _08183_ (.A1_N(_02658_),
    .A2_N(_02659_),
    .B1(_02656_),
    .B2(_01911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[5] ));
 sky130_fd_sc_hd__o22a_1 _08184_ (.A1(_02595_),
    .A2(_02606_),
    .B1(_02609_),
    .B2(_02640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02660_));
 sky130_fd_sc_hd__a31o_1 _08185_ (.A1(_02653_),
    .A2(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .A3(_02621_),
    .B1(_02637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02661_));
 sky130_fd_sc_hd__and3_1 _08186_ (.A(_02583_),
    .B(_02660_),
    .C(_02661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02662_));
 sky130_fd_sc_hd__and2_1 _08187_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[6] ),
    .B(_02662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02663_));
 sky130_fd_sc_hd__nor2_1 _08188_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[6] ),
    .B(_02662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02664_));
 sky130_fd_sc_hd__or2_1 _08189_ (.A(_02663_),
    .B(_02664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02665_));
 sky130_fd_sc_hd__a22o_1 _08190_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[4] ),
    .A2(_02642_),
    .B1(_02656_),
    .B2(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02666_));
 sky130_fd_sc_hd__o21ai_1 _08191_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[5] ),
    .A2(_02656_),
    .B1(_02666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02667_));
 sky130_fd_sc_hd__o41a_2 _08192_ (.A1(_02628_),
    .A2(_02645_),
    .A3(_02646_),
    .A4(_02657_),
    .B1(_02667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02668_));
 sky130_fd_sc_hd__xor2_1 _08193_ (.A(_02665_),
    .B(_02668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02669_));
 sky130_fd_sc_hd__mux2_1 _08194_ (.A0(_02662_),
    .A1(_02669_),
    .S(_02618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02670_));
 sky130_fd_sc_hd__clkbuf_1 _08195_ (.A(_02670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[6] ));
 sky130_fd_sc_hd__o22a_1 _08196_ (.A1(_02595_),
    .A2(_02620_),
    .B1(_02625_),
    .B2(_02640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02671_));
 sky130_fd_sc_hd__clkbuf_4 _08197_ (.A(_02621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02672_));
 sky130_fd_sc_hd__a31o_1 _08198_ (.A1(_02653_),
    .A2(_02672_),
    .A3(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .B1(_02637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02673_));
 sky130_fd_sc_hd__and3_1 _08199_ (.A(_02583_),
    .B(_02671_),
    .C(_02673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02674_));
 sky130_fd_sc_hd__and2_1 _08200_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[7] ),
    .B(_02674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02675_));
 sky130_fd_sc_hd__nor2_1 _08201_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[7] ),
    .B(_02674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02676_));
 sky130_fd_sc_hd__or2_1 _08202_ (.A(_02675_),
    .B(_02676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02677_));
 sky130_fd_sc_hd__o21bai_1 _08203_ (.A1(_02665_),
    .A2(_02668_),
    .B1_N(_02663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02678_));
 sky130_fd_sc_hd__xnor2_1 _08204_ (.A(_02677_),
    .B(_02678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02679_));
 sky130_fd_sc_hd__mux2_1 _08205_ (.A0(_02674_),
    .A1(_02679_),
    .S(_02618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02680_));
 sky130_fd_sc_hd__clkbuf_1 _08206_ (.A(_02680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[7] ));
 sky130_fd_sc_hd__and3_1 _08207_ (.A(_02654_),
    .B(_02584_),
    .C(_02588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02681_));
 sky130_fd_sc_hd__nor2_1 _08208_ (.A(_02586_),
    .B(\sa_inst.sak._13_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02682_));
 sky130_fd_sc_hd__and3_1 _08209_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[8] ),
    .B(_02588_),
    .C(_02682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02683_));
 sky130_fd_sc_hd__nor2_1 _08210_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[8] ),
    .B(_02681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02684_));
 sky130_fd_sc_hd__or2_1 _08211_ (.A(_02683_),
    .B(_02684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02685_));
 sky130_fd_sc_hd__o21bai_1 _08212_ (.A1(_02663_),
    .A2(_02675_),
    .B1_N(_02676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02686_));
 sky130_fd_sc_hd__o31ai_2 _08213_ (.A1(_02665_),
    .A2(_02668_),
    .A3(_02677_),
    .B1(_02686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02687_));
 sky130_fd_sc_hd__xnor2_1 _08214_ (.A(_02685_),
    .B(_02687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02688_));
 sky130_fd_sc_hd__mux2_1 _08215_ (.A0(_02681_),
    .A1(_02688_),
    .S(_02618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02689_));
 sky130_fd_sc_hd__clkbuf_1 _08216_ (.A(_02689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[8] ));
 sky130_fd_sc_hd__buf_2 _08217_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02690_));
 sky130_fd_sc_hd__clkbuf_4 _08218_ (.A(_02690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02691_));
 sky130_fd_sc_hd__and3_1 _08219_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[9] ),
    .B(_02598_),
    .C(_02682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02692_));
 sky130_fd_sc_hd__and3_1 _08220_ (.A(_02654_),
    .B(_02584_),
    .C(_02598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02693_));
 sky130_fd_sc_hd__nor2_1 _08221_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[9] ),
    .B(_02693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02694_));
 sky130_fd_sc_hd__or2_1 _08222_ (.A(_02692_),
    .B(_02694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02695_));
 sky130_fd_sc_hd__inv_2 _08223_ (.A(_02685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02696_));
 sky130_fd_sc_hd__a21oi_1 _08224_ (.A1(_02696_),
    .A2(_02687_),
    .B1(_02683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02697_));
 sky130_fd_sc_hd__xnor2_1 _08225_ (.A(_02695_),
    .B(_02697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02698_));
 sky130_fd_sc_hd__nor2_1 _08226_ (.A(_01978_),
    .B(_02693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02699_));
 sky130_fd_sc_hd__a21oi_1 _08227_ (.A1(_02691_),
    .A2(_02698_),
    .B1(_02699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[9] ));
 sky130_fd_sc_hd__mux2_1 _08228_ (.A0(_02606_),
    .A1(_02607_),
    .S(_02610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02700_));
 sky130_fd_sc_hd__and2_1 _08229_ (.A(_02700_),
    .B(_02682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02701_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08230_ (.A(_02682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02702_));
 sky130_fd_sc_hd__and3_1 _08231_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[10] ),
    .B(_02700_),
    .C(_02702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02703_));
 sky130_fd_sc_hd__nor2_1 _08232_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[10] ),
    .B(_02701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02704_));
 sky130_fd_sc_hd__or2_1 _08233_ (.A(_02703_),
    .B(_02704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02705_));
 sky130_fd_sc_hd__inv_2 _08234_ (.A(_02694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02706_));
 sky130_fd_sc_hd__a211o_1 _08235_ (.A1(_02696_),
    .A2(_02687_),
    .B1(_02692_),
    .C1(_02683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02707_));
 sky130_fd_sc_hd__and2_1 _08236_ (.A(_02706_),
    .B(_02707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02708_));
 sky130_fd_sc_hd__xnor2_1 _08237_ (.A(_02705_),
    .B(_02708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02709_));
 sky130_fd_sc_hd__buf_2 _08238_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02710_));
 sky130_fd_sc_hd__mux2_1 _08239_ (.A0(_02701_),
    .A1(_02709_),
    .S(_02710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02711_));
 sky130_fd_sc_hd__clkbuf_1 _08240_ (.A(_02711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[10] ));
 sky130_fd_sc_hd__o211a_1 _08241_ (.A1(_02610_),
    .A2(_02620_),
    .B1(_02623_),
    .C1(_02702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02712_));
 sky130_fd_sc_hd__and2_1 _08242_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[11] ),
    .B(_02712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02713_));
 sky130_fd_sc_hd__or2_1 _08243_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[11] ),
    .B(_02712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02714_));
 sky130_fd_sc_hd__or2b_1 _08244_ (.A(_02713_),
    .B_N(_02714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02715_));
 sky130_fd_sc_hd__inv_2 _08245_ (.A(_02704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02716_));
 sky130_fd_sc_hd__a31o_1 _08246_ (.A1(_02706_),
    .A2(_02716_),
    .A3(_02707_),
    .B1(_02703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02717_));
 sky130_fd_sc_hd__xnor2_1 _08247_ (.A(_02715_),
    .B(_02717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02718_));
 sky130_fd_sc_hd__mux2_1 _08248_ (.A0(_02712_),
    .A1(_02718_),
    .S(_02710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02719_));
 sky130_fd_sc_hd__clkbuf_1 _08249_ (.A(_02719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[11] ));
 sky130_fd_sc_hd__and3_1 _08250_ (.A(_02653_),
    .B(_02636_),
    .C(_02682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02720_));
 sky130_fd_sc_hd__and2_1 _08251_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[12] ),
    .B(_02720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02721_));
 sky130_fd_sc_hd__nor2_1 _08252_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[12] ),
    .B(_02720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02722_));
 sky130_fd_sc_hd__or2_1 _08253_ (.A(_02721_),
    .B(_02722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02723_));
 sky130_fd_sc_hd__inv_2 _08254_ (.A(_02723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02724_));
 sky130_fd_sc_hd__a311o_1 _08255_ (.A1(_02706_),
    .A2(_02716_),
    .A3(_02707_),
    .B1(_02713_),
    .C1(_02703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02725_));
 sky130_fd_sc_hd__nand2_1 _08256_ (.A(_02714_),
    .B(_02725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02726_));
 sky130_fd_sc_hd__xnor2_1 _08257_ (.A(_02724_),
    .B(_02726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02727_));
 sky130_fd_sc_hd__mux2_1 _08258_ (.A0(_02720_),
    .A1(_02727_),
    .S(_02710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02728_));
 sky130_fd_sc_hd__clkbuf_1 _08259_ (.A(_02728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[12] ));
 sky130_fd_sc_hd__buf_2 _08260_ (.A(_02690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02729_));
 sky130_fd_sc_hd__clkbuf_2 _08261_ (.A(_02653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02730_));
 sky130_fd_sc_hd__and3_1 _08262_ (.A(_02730_),
    .B(_02651_),
    .C(_02702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02731_));
 sky130_fd_sc_hd__and2_1 _08263_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[13] ),
    .B(_02731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02732_));
 sky130_fd_sc_hd__nor2_1 _08264_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[13] ),
    .B(_02731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02733_));
 sky130_fd_sc_hd__nor2_1 _08265_ (.A(_02732_),
    .B(_02733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02734_));
 sky130_fd_sc_hd__a31o_1 _08266_ (.A1(_02714_),
    .A2(_02724_),
    .A3(_02725_),
    .B1(_02721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02735_));
 sky130_fd_sc_hd__xnor2_1 _08267_ (.A(_02734_),
    .B(_02735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02736_));
 sky130_fd_sc_hd__nor2_1 _08268_ (.A(_01978_),
    .B(_02731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02737_));
 sky130_fd_sc_hd__a21oi_1 _08269_ (.A1(_02729_),
    .A2(_02736_),
    .B1(_02737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[13] ));
 sky130_fd_sc_hd__and3_1 _08270_ (.A(_02730_),
    .B(_02607_),
    .C(_02702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02738_));
 sky130_fd_sc_hd__and2_1 _08271_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[14] ),
    .B(_02738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02739_));
 sky130_fd_sc_hd__nor2_1 _08272_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[14] ),
    .B(_02738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02740_));
 sky130_fd_sc_hd__or2_1 _08273_ (.A(_02739_),
    .B(_02740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02741_));
 sky130_fd_sc_hd__o21ba_1 _08274_ (.A1(_02721_),
    .A2(_02732_),
    .B1_N(_02733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02742_));
 sky130_fd_sc_hd__a41o_1 _08275_ (.A1(_02714_),
    .A2(_02724_),
    .A3(_02725_),
    .A4(_02734_),
    .B1(_02742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02743_));
 sky130_fd_sc_hd__xnor2_1 _08276_ (.A(_02741_),
    .B(_02743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02744_));
 sky130_fd_sc_hd__mux2_1 _08277_ (.A0(_02738_),
    .A1(_02744_),
    .S(_02710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02745_));
 sky130_fd_sc_hd__clkbuf_1 _08278_ (.A(_02745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[14] ));
 sky130_fd_sc_hd__and4_1 _08279_ (.A(_02730_),
    .B(_02672_),
    .C(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .D(_02702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02746_));
 sky130_fd_sc_hd__and2_1 _08280_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[15] ),
    .B(_02746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02747_));
 sky130_fd_sc_hd__nor2_1 _08281_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[15] ),
    .B(_02746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02748_));
 sky130_fd_sc_hd__nor2_1 _08282_ (.A(_02747_),
    .B(_02748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02749_));
 sky130_fd_sc_hd__inv_2 _08283_ (.A(_02741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02750_));
 sky130_fd_sc_hd__a21oi_1 _08284_ (.A1(_02750_),
    .A2(_02743_),
    .B1(_02739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02751_));
 sky130_fd_sc_hd__xnor2_1 _08285_ (.A(_02749_),
    .B(_02751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02752_));
 sky130_fd_sc_hd__mux2_1 _08286_ (.A0(_02746_),
    .A1(_02752_),
    .S(_02710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02753_));
 sky130_fd_sc_hd__clkbuf_1 _08287_ (.A(_02753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[15] ));
 sky130_fd_sc_hd__o21ba_1 _08288_ (.A1(_02739_),
    .A2(_02747_),
    .B1_N(_02748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02754_));
 sky130_fd_sc_hd__a31o_1 _08289_ (.A1(_02750_),
    .A2(_02743_),
    .A3(_02749_),
    .B1(_02754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02755_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08290_ (.A(_02755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02756_));
 sky130_fd_sc_hd__a21oi_1 _08291_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[16] ),
    .A2(_02756_),
    .B1(_02635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02757_));
 sky130_fd_sc_hd__o21a_1 _08292_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[16] ),
    .A2(_02756_),
    .B1(_02757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[16] ));
 sky130_fd_sc_hd__and2_1 _08293_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[16] ),
    .B(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02758_));
 sky130_fd_sc_hd__and2_1 _08294_ (.A(_02756_),
    .B(_02758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02759_));
 sky130_fd_sc_hd__a21o_1 _08295_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[16] ),
    .A2(_02756_),
    .B1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02760_));
 sky130_fd_sc_hd__and3b_1 _08296_ (.A_N(_02759_),
    .B(_01828_),
    .C(_02760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02761_));
 sky130_fd_sc_hd__clkbuf_1 _08297_ (.A(_02761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[17] ));
 sky130_fd_sc_hd__clkbuf_2 _08298_ (.A(_02690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02762_));
 sky130_fd_sc_hd__o21ai_1 _08299_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[18] ),
    .A2(_02759_),
    .B1(_02762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02763_));
 sky130_fd_sc_hd__a21oi_1 _08300_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[18] ),
    .A2(_02759_),
    .B1(_02763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[18] ));
 sky130_fd_sc_hd__and4_1 _08301_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[18] ),
    .B(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[19] ),
    .C(_02755_),
    .D(_02758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02764_));
 sky130_fd_sc_hd__clkbuf_1 _08302_ (.A(_02764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02765_));
 sky130_fd_sc_hd__buf_4 _08303_ (.A(_01825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02766_));
 sky130_fd_sc_hd__a31o_1 _08304_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[18] ),
    .A2(_02756_),
    .A3(_02758_),
    .B1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02767_));
 sky130_fd_sc_hd__and3b_1 _08305_ (.A_N(_02765_),
    .B(_02766_),
    .C(_02767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02768_));
 sky130_fd_sc_hd__clkbuf_1 _08306_ (.A(_02768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[19] ));
 sky130_fd_sc_hd__and2_1 _08307_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[20] ),
    .B(_02765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02769_));
 sky130_fd_sc_hd__o21ai_1 _08308_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[20] ),
    .A2(_02765_),
    .B1(_02729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02770_));
 sky130_fd_sc_hd__nor2_1 _08309_ (.A(_02769_),
    .B(_02770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[20] ));
 sky130_fd_sc_hd__and2_1 _08310_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[20] ),
    .B(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02771_));
 sky130_fd_sc_hd__and2_1 _08311_ (.A(_02765_),
    .B(_02771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02772_));
 sky130_fd_sc_hd__inv_2 _08312_ (.A(_02772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02773_));
 sky130_fd_sc_hd__o211a_1 _08313_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[21] ),
    .A2(_02769_),
    .B1(_02773_),
    .C1(_01829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[21] ));
 sky130_fd_sc_hd__and3_1 _08314_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[22] ),
    .B(_02765_),
    .C(_02771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02774_));
 sky130_fd_sc_hd__o21ai_1 _08315_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[22] ),
    .A2(_02772_),
    .B1(_02729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02775_));
 sky130_fd_sc_hd__nor2_1 _08316_ (.A(_02774_),
    .B(_02775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[22] ));
 sky130_fd_sc_hd__and4_1 _08317_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[22] ),
    .B(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[23] ),
    .C(_02764_),
    .D(_02771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02776_));
 sky130_fd_sc_hd__o21ai_1 _08318_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[23] ),
    .A2(_02774_),
    .B1(_02729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02777_));
 sky130_fd_sc_hd__nor2_1 _08319_ (.A(_02776_),
    .B(_02777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[23] ));
 sky130_fd_sc_hd__and2_1 _08320_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[24] ),
    .B(_02776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02778_));
 sky130_fd_sc_hd__o21ai_1 _08321_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[24] ),
    .A2(_02776_),
    .B1(_02762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02779_));
 sky130_fd_sc_hd__nor2_1 _08322_ (.A(_02778_),
    .B(_02779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[24] ));
 sky130_fd_sc_hd__o21ai_1 _08323_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[25] ),
    .A2(_02778_),
    .B1(_02762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02780_));
 sky130_fd_sc_hd__a21oi_1 _08324_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[25] ),
    .A2(_02778_),
    .B1(_02780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[25] ));
 sky130_fd_sc_hd__and4_1 _08325_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[24] ),
    .B(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[25] ),
    .C(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[26] ),
    .D(_02776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02781_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08326_ (.A(_02781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02782_));
 sky130_fd_sc_hd__a31o_1 _08327_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[24] ),
    .A2(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[25] ),
    .A3(_02776_),
    .B1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02783_));
 sky130_fd_sc_hd__and3b_1 _08328_ (.A_N(_02782_),
    .B(_02766_),
    .C(_02783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02784_));
 sky130_fd_sc_hd__clkbuf_1 _08329_ (.A(_02784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[26] ));
 sky130_fd_sc_hd__clkbuf_1 _08330_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02785_));
 sky130_fd_sc_hd__and2_1 _08331_ (.A(_02785_),
    .B(_02782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02786_));
 sky130_fd_sc_hd__o21ai_1 _08332_ (.A1(_02785_),
    .A2(_02782_),
    .B1(_02762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02787_));
 sky130_fd_sc_hd__nor2_1 _08333_ (.A(_02786_),
    .B(_02787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[27] ));
 sky130_fd_sc_hd__o21ai_1 _08334_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[28] ),
    .A2(_02786_),
    .B1(_02762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02788_));
 sky130_fd_sc_hd__a21oi_1 _08335_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[28] ),
    .A2(_02786_),
    .B1(_02788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[28] ));
 sky130_fd_sc_hd__and2_1 _08336_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[28] ),
    .B(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02789_));
 sky130_fd_sc_hd__a31o_1 _08337_ (.A1(_02785_),
    .A2(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[28] ),
    .A3(_02782_),
    .B1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02790_));
 sky130_fd_sc_hd__nand2_1 _08338_ (.A(_02729_),
    .B(_02790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02791_));
 sky130_fd_sc_hd__a21oi_1 _08339_ (.A1(_02786_),
    .A2(_02789_),
    .B1(_02791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[29] ));
 sky130_fd_sc_hd__and4_1 _08340_ (.A(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[27] ),
    .B(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[30] ),
    .C(_02781_),
    .D(_02789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02792_));
 sky130_fd_sc_hd__a31o_1 _08341_ (.A1(_02785_),
    .A2(_02782_),
    .A3(_02789_),
    .B1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02793_));
 sky130_fd_sc_hd__and3b_1 _08342_ (.A_N(_02792_),
    .B(_02766_),
    .C(_02793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02794_));
 sky130_fd_sc_hd__clkbuf_1 _08343_ (.A(_02794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[30] ));
 sky130_fd_sc_hd__a21oi_1 _08344_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[31] ),
    .A2(_02792_),
    .B1(_02635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02795_));
 sky130_fd_sc_hd__o21a_1 _08345_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[31] ),
    .A2(_02792_),
    .B1(_02795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[31] ));
 sky130_fd_sc_hd__buf_4 _08346_ (.A(\sa_inst.sak._21_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02796_));
 sky130_fd_sc_hd__buf_2 _08347_ (.A(_02796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02797_));
 sky130_fd_sc_hd__mux2_1 _08348_ (.A0(\sa_inst.sak._01_[0] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[0] ),
    .S(_02797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02798_));
 sky130_fd_sc_hd__clkbuf_1 _08349_ (.A(_02798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ));
 sky130_fd_sc_hd__mux2_1 _08350_ (.A0(\sa_inst.sak._01_[1] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[1] ),
    .S(_02797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02799_));
 sky130_fd_sc_hd__clkbuf_1 _08351_ (.A(_02799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ));
 sky130_fd_sc_hd__clkbuf_4 _08352_ (.A(\sa_inst.sak._21_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02800_));
 sky130_fd_sc_hd__clkbuf_2 _08353_ (.A(_02800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02801_));
 sky130_fd_sc_hd__mux2_1 _08354_ (.A0(\sa_inst.sak._01_[2] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[2] ),
    .S(_02801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02802_));
 sky130_fd_sc_hd__clkbuf_1 _08355_ (.A(_02802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ));
 sky130_fd_sc_hd__mux2_1 _08356_ (.A0(\sa_inst.sak._01_[3] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[3] ),
    .S(_02801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02803_));
 sky130_fd_sc_hd__clkbuf_1 _08357_ (.A(_02803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ));
 sky130_fd_sc_hd__mux2_1 _08358_ (.A0(\sa_inst.sak._01_[4] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[4] ),
    .S(_02801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02804_));
 sky130_fd_sc_hd__clkbuf_1 _08359_ (.A(_02804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ));
 sky130_fd_sc_hd__mux2_1 _08360_ (.A0(\sa_inst.sak._01_[5] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[5] ),
    .S(_02801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02805_));
 sky130_fd_sc_hd__clkbuf_1 _08361_ (.A(_02805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ));
 sky130_fd_sc_hd__mux2_1 _08362_ (.A0(\sa_inst.sak._01_[6] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[6] ),
    .S(_02801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02806_));
 sky130_fd_sc_hd__clkbuf_1 _08363_ (.A(_02806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ));
 sky130_fd_sc_hd__clkbuf_2 _08364_ (.A(_02800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02807_));
 sky130_fd_sc_hd__mux2_1 _08365_ (.A0(\sa_inst.sak._01_[7] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[7] ),
    .S(_02807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02808_));
 sky130_fd_sc_hd__clkbuf_1 _08366_ (.A(_02808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ));
 sky130_fd_sc_hd__mux2_1 _08367_ (.A0(\sa_inst.sak._01_[8] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[8] ),
    .S(_02807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02809_));
 sky130_fd_sc_hd__clkbuf_1 _08368_ (.A(_02809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ));
 sky130_fd_sc_hd__mux2_1 _08369_ (.A0(\sa_inst.sak._01_[9] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[9] ),
    .S(_02807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02810_));
 sky130_fd_sc_hd__clkbuf_1 _08370_ (.A(_02810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ));
 sky130_fd_sc_hd__mux2_1 _08371_ (.A0(\sa_inst.sak._01_[10] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[10] ),
    .S(_02807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02811_));
 sky130_fd_sc_hd__clkbuf_1 _08372_ (.A(_02811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ));
 sky130_fd_sc_hd__mux2_1 _08373_ (.A0(\sa_inst.sak._01_[11] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[11] ),
    .S(_02807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02812_));
 sky130_fd_sc_hd__clkbuf_1 _08374_ (.A(_02812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ));
 sky130_fd_sc_hd__buf_2 _08375_ (.A(_02800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02813_));
 sky130_fd_sc_hd__mux2_1 _08376_ (.A0(\sa_inst.sak._01_[12] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[12] ),
    .S(_02813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02814_));
 sky130_fd_sc_hd__clkbuf_1 _08377_ (.A(_02814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ));
 sky130_fd_sc_hd__mux2_1 _08378_ (.A0(\sa_inst.sak._01_[13] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[13] ),
    .S(_02813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02815_));
 sky130_fd_sc_hd__clkbuf_1 _08379_ (.A(_02815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ));
 sky130_fd_sc_hd__mux2_1 _08380_ (.A0(\sa_inst.sak._01_[14] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[14] ),
    .S(_02813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02816_));
 sky130_fd_sc_hd__clkbuf_1 _08381_ (.A(_02816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ));
 sky130_fd_sc_hd__mux2_1 _08382_ (.A0(\sa_inst.sak._01_[15] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[15] ),
    .S(_02813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02817_));
 sky130_fd_sc_hd__clkbuf_1 _08383_ (.A(_02817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ));
 sky130_fd_sc_hd__mux2_1 _08384_ (.A0(\sa_inst.sak._01_[16] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[16] ),
    .S(_02813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02818_));
 sky130_fd_sc_hd__clkbuf_1 _08385_ (.A(_02818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ));
 sky130_fd_sc_hd__clkbuf_2 _08386_ (.A(_02800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02819_));
 sky130_fd_sc_hd__mux2_1 _08387_ (.A0(\sa_inst.sak._01_[17] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[17] ),
    .S(_02819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02820_));
 sky130_fd_sc_hd__clkbuf_1 _08388_ (.A(_02820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ));
 sky130_fd_sc_hd__mux2_1 _08389_ (.A0(\sa_inst.sak._01_[18] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[18] ),
    .S(_02819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02821_));
 sky130_fd_sc_hd__clkbuf_1 _08390_ (.A(_02821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ));
 sky130_fd_sc_hd__mux2_1 _08391_ (.A0(\sa_inst.sak._01_[19] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[19] ),
    .S(_02819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02822_));
 sky130_fd_sc_hd__clkbuf_1 _08392_ (.A(_02822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ));
 sky130_fd_sc_hd__mux2_1 _08393_ (.A0(\sa_inst.sak._01_[20] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[20] ),
    .S(_02819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02823_));
 sky130_fd_sc_hd__clkbuf_1 _08394_ (.A(_02823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ));
 sky130_fd_sc_hd__mux2_1 _08395_ (.A0(\sa_inst.sak._01_[21] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[21] ),
    .S(_02819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02824_));
 sky130_fd_sc_hd__clkbuf_1 _08396_ (.A(_02824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ));
 sky130_fd_sc_hd__clkbuf_2 _08397_ (.A(_02800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02825_));
 sky130_fd_sc_hd__mux2_1 _08398_ (.A0(\sa_inst.sak._01_[22] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[22] ),
    .S(_02825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02826_));
 sky130_fd_sc_hd__clkbuf_1 _08399_ (.A(_02826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ));
 sky130_fd_sc_hd__mux2_1 _08400_ (.A0(\sa_inst.sak._01_[23] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[23] ),
    .S(_02825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02827_));
 sky130_fd_sc_hd__clkbuf_1 _08401_ (.A(_02827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ));
 sky130_fd_sc_hd__mux2_1 _08402_ (.A0(\sa_inst.sak._01_[24] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[24] ),
    .S(_02825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02828_));
 sky130_fd_sc_hd__clkbuf_1 _08403_ (.A(_02828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ));
 sky130_fd_sc_hd__mux2_1 _08404_ (.A0(\sa_inst.sak._01_[25] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[25] ),
    .S(_02825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02829_));
 sky130_fd_sc_hd__clkbuf_1 _08405_ (.A(_02829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ));
 sky130_fd_sc_hd__mux2_1 _08406_ (.A0(\sa_inst.sak._01_[26] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[26] ),
    .S(_02825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02830_));
 sky130_fd_sc_hd__clkbuf_1 _08407_ (.A(_02830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ));
 sky130_fd_sc_hd__clkbuf_4 _08408_ (.A(\sa_inst.sak._21_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02831_));
 sky130_fd_sc_hd__clkbuf_2 _08409_ (.A(_02831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02832_));
 sky130_fd_sc_hd__mux2_1 _08410_ (.A0(\sa_inst.sak._01_[27] ),
    .A1(_02785_),
    .S(_02832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02833_));
 sky130_fd_sc_hd__clkbuf_1 _08411_ (.A(_02833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ));
 sky130_fd_sc_hd__mux2_1 _08412_ (.A0(\sa_inst.sak._01_[28] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[28] ),
    .S(_02832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02834_));
 sky130_fd_sc_hd__clkbuf_1 _08413_ (.A(_02834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ));
 sky130_fd_sc_hd__mux2_1 _08414_ (.A0(\sa_inst.sak._01_[29] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[29] ),
    .S(_02832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02835_));
 sky130_fd_sc_hd__clkbuf_1 _08415_ (.A(_02835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ));
 sky130_fd_sc_hd__mux2_1 _08416_ (.A0(\sa_inst.sak._01_[30] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[30] ),
    .S(_02832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02836_));
 sky130_fd_sc_hd__clkbuf_1 _08417_ (.A(_02836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ));
 sky130_fd_sc_hd__mux2_1 _08418_ (.A0(\sa_inst.sak._01_[31] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[31] ),
    .S(_02832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02837_));
 sky130_fd_sc_hd__clkbuf_1 _08419_ (.A(_02837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ));
 sky130_fd_sc_hd__buf_2 _08420_ (.A(_02831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02838_));
 sky130_fd_sc_hd__mux2_1 _08421_ (.A0(\sa_inst.sak._01_[32] ),
    .A1(\sa_inst.sak.rows:2.cols:2.pe_ij._02_ ),
    .S(_02838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02839_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08422_ (.A(_02839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ));
 sky130_fd_sc_hd__xor2_2 _08423_ (.A(\sa_inst.sak._03_[10] ),
    .B(\sa_inst.sak._13_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02840_));
 sky130_fd_sc_hd__clkbuf_2 _08424_ (.A(_02840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02841_));
 sky130_fd_sc_hd__clkbuf_2 _08425_ (.A(_02841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._01_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08426_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._00_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02842_));
 sky130_fd_sc_hd__clkbuf_4 _08427_ (.A(_02842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02843_));
 sky130_fd_sc_hd__inv_2 _08428_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02844_));
 sky130_fd_sc_hd__clkbuf_2 _08429_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02845_));
 sky130_fd_sc_hd__mux2_1 _08430_ (.A0(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[1] ),
    .S(_02845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02846_));
 sky130_fd_sc_hd__and2b_1 _08431_ (.A_N(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._22_ ),
    .B(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02847_));
 sky130_fd_sc_hd__clkbuf_2 _08432_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02848_));
 sky130_fd_sc_hd__mux4_1 _08433_ (.A0(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .A2(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .A3(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .S0(_02848_),
    .S1(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02849_));
 sky130_fd_sc_hd__nor2_2 _08434_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._22_ ),
    .B(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02850_));
 sky130_fd_sc_hd__a32o_2 _08435_ (.A1(_02844_),
    .A2(_02846_),
    .A3(_02847_),
    .B1(_02849_),
    .B2(_02850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02851_));
 sky130_fd_sc_hd__xor2_4 _08436_ (.A(_02843_),
    .B(_02851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02852_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08437_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02853_));
 sky130_fd_sc_hd__buf_2 _08438_ (.A(_02853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02854_));
 sky130_fd_sc_hd__nand2_1 _08439_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[0] ),
    .B(_02854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02855_));
 sky130_fd_sc_hd__xnor2_1 _08440_ (.A(_02852_),
    .B(_02855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[0] ));
 sky130_fd_sc_hd__inv_2 _08441_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._22_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02856_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08442_ (.A(_02856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02857_));
 sky130_fd_sc_hd__mux2_1 _08443_ (.A0(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .S(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02858_));
 sky130_fd_sc_hd__mux2_1 _08444_ (.A0(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .S(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02859_));
 sky130_fd_sc_hd__mux2_1 _08445_ (.A0(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[2] ),
    .S(_02848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02860_));
 sky130_fd_sc_hd__and2b_1 _08446_ (.A_N(_02845_),
    .B(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02861_));
 sky130_fd_sc_hd__clkbuf_2 _08447_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02862_));
 sky130_fd_sc_hd__clkbuf_2 _08448_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02863_));
 sky130_fd_sc_hd__mux4_2 _08449_ (.A0(_02858_),
    .A1(_02859_),
    .A2(_02860_),
    .A3(_02861_),
    .S0(_02862_),
    .S1(_02863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02864_));
 sky130_fd_sc_hd__nand4_2 _08450_ (.A(_02857_),
    .B(_02843_),
    .C(_02851_),
    .D(_02864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02865_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08451_ (.A(_02865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02866_));
 sky130_fd_sc_hd__clkbuf_2 _08452_ (.A(_02857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02867_));
 sky130_fd_sc_hd__a22o_1 _08453_ (.A1(_02843_),
    .A2(_02851_),
    .B1(_02864_),
    .B2(_02867_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02868_));
 sky130_fd_sc_hd__and2_1 _08454_ (.A(_02866_),
    .B(_02868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02869_));
 sky130_fd_sc_hd__and3_1 _08455_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[1] ),
    .B(_02865_),
    .C(_02868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02870_));
 sky130_fd_sc_hd__a21oi_1 _08456_ (.A1(_02866_),
    .A2(_02868_),
    .B1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02871_));
 sky130_fd_sc_hd__or2_1 _08457_ (.A(_02870_),
    .B(_02871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02872_));
 sky130_fd_sc_hd__nand2_1 _08458_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[0] ),
    .B(_02852_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02873_));
 sky130_fd_sc_hd__xor2_1 _08459_ (.A(_02872_),
    .B(_02873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02874_));
 sky130_fd_sc_hd__buf_2 _08460_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02875_));
 sky130_fd_sc_hd__mux2_1 _08461_ (.A0(_02869_),
    .A1(_02874_),
    .S(_02875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02876_));
 sky130_fd_sc_hd__clkbuf_1 _08462_ (.A(_02876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[1] ));
 sky130_fd_sc_hd__clkbuf_4 _08463_ (.A(_02853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02877_));
 sky130_fd_sc_hd__buf_2 _08464_ (.A(_02877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02878_));
 sky130_fd_sc_hd__o21ba_1 _08465_ (.A1(_02871_),
    .A2(_02873_),
    .B1_N(_02870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02879_));
 sky130_fd_sc_hd__mux2_1 _08466_ (.A0(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._00_ ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .S(_02848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02880_));
 sky130_fd_sc_hd__mux2_1 _08467_ (.A0(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .S(_02848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02881_));
 sky130_fd_sc_hd__clkbuf_2 _08468_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02882_));
 sky130_fd_sc_hd__mux2_1 _08469_ (.A0(_02880_),
    .A1(_02881_),
    .S(_02882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02883_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08470_ (.A(_02844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02884_));
 sky130_fd_sc_hd__mux2_1 _08471_ (.A0(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ),
    .S(_02845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02885_));
 sky130_fd_sc_hd__clkbuf_2 _08472_ (.A(_02848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02886_));
 sky130_fd_sc_hd__and3b_1 _08473_ (.A_N(_02886_),
    .B(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[1] ),
    .C(_02862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02887_));
 sky130_fd_sc_hd__a21o_1 _08474_ (.A1(_02884_),
    .A2(_02885_),
    .B1(_02887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02888_));
 sky130_fd_sc_hd__a22oi_4 _08475_ (.A1(_02850_),
    .A2(_02883_),
    .B1(_02888_),
    .B2(_02847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02889_));
 sky130_fd_sc_hd__xor2_1 _08476_ (.A(_02865_),
    .B(_02889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02890_));
 sky130_fd_sc_hd__nor2_1 _08477_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[2] ),
    .B(_02890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02891_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08478_ (.A(_02890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02892_));
 sky130_fd_sc_hd__nand2_1 _08479_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[2] ),
    .B(_02892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02893_));
 sky130_fd_sc_hd__and2b_1 _08480_ (.A_N(_02891_),
    .B(_02893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02894_));
 sky130_fd_sc_hd__xnor2_1 _08481_ (.A(_02879_),
    .B(_02894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02895_));
 sky130_fd_sc_hd__inv_2 _08482_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02896_));
 sky130_fd_sc_hd__buf_2 _08483_ (.A(_02896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02897_));
 sky130_fd_sc_hd__clkbuf_4 _08484_ (.A(_02897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02898_));
 sky130_fd_sc_hd__and2_1 _08485_ (.A(_02898_),
    .B(_02892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02899_));
 sky130_fd_sc_hd__a21o_1 _08486_ (.A1(_02878_),
    .A2(_02895_),
    .B1(_02899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[2] ));
 sky130_fd_sc_hd__mux4_2 _08487_ (.A0(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._00_ ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .A2(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .A3(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .S0(_02862_),
    .S1(_02886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02900_));
 sky130_fd_sc_hd__mux4_1 _08488_ (.A0(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[2] ),
    .A2(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ),
    .A3(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[0] ),
    .S0(_02862_),
    .S1(_02886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02901_));
 sky130_fd_sc_hd__a22o_1 _08489_ (.A1(_02850_),
    .A2(_02900_),
    .B1(_02901_),
    .B2(_02847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02902_));
 sky130_fd_sc_hd__nor3b_1 _08490_ (.A(_02865_),
    .B(_02889_),
    .C_N(_02902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02903_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08491_ (.A(_02903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02904_));
 sky130_fd_sc_hd__o21bai_1 _08492_ (.A1(_02866_),
    .A2(_02889_),
    .B1_N(_02902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02905_));
 sky130_fd_sc_hd__and2b_1 _08493_ (.A_N(_02904_),
    .B(_02905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02906_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08494_ (.A(_02906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02907_));
 sky130_fd_sc_hd__nor2_1 _08495_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[3] ),
    .B(_02906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02908_));
 sky130_fd_sc_hd__buf_2 _08496_ (.A(_02903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02909_));
 sky130_fd_sc_hd__nand3b_1 _08497_ (.A_N(_02909_),
    .B(_02905_),
    .C(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02910_));
 sky130_fd_sc_hd__or2b_1 _08498_ (.A(_02908_),
    .B_N(_02910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02911_));
 sky130_fd_sc_hd__o21a_1 _08499_ (.A1(_02879_),
    .A2(_02891_),
    .B1(_02893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02912_));
 sky130_fd_sc_hd__xor2_1 _08500_ (.A(_02911_),
    .B(_02912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02913_));
 sky130_fd_sc_hd__buf_2 _08501_ (.A(_02853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02914_));
 sky130_fd_sc_hd__mux2_1 _08502_ (.A0(_02907_),
    .A1(_02913_),
    .S(_02914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02915_));
 sky130_fd_sc_hd__clkbuf_1 _08503_ (.A(_02915_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[3] ));
 sky130_fd_sc_hd__clkbuf_4 _08504_ (.A(_02854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02916_));
 sky130_fd_sc_hd__mux2_1 _08505_ (.A0(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .S(_02845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02917_));
 sky130_fd_sc_hd__mux2_1 _08506_ (.A0(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .S(_02845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02918_));
 sky130_fd_sc_hd__mux4_1 _08507_ (.A0(_02842_),
    .A1(_02917_),
    .A2(_02918_),
    .A3(_02846_),
    .S0(_02882_),
    .S1(_02863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02919_));
 sky130_fd_sc_hd__and2_1 _08508_ (.A(_02867_),
    .B(_02919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02920_));
 sky130_fd_sc_hd__xor2_4 _08509_ (.A(_02909_),
    .B(_02920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02921_));
 sky130_fd_sc_hd__xnor2_1 _08510_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[4] ),
    .B(_02921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02922_));
 sky130_fd_sc_hd__o211a_1 _08511_ (.A1(_02879_),
    .A2(_02891_),
    .B1(_02893_),
    .C1(_02910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02923_));
 sky130_fd_sc_hd__or3_1 _08512_ (.A(_02908_),
    .B(_02922_),
    .C(_02923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02924_));
 sky130_fd_sc_hd__o21ai_1 _08513_ (.A1(_02908_),
    .A2(_02923_),
    .B1(_02922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02925_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08514_ (.A(_02897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02926_));
 sky130_fd_sc_hd__and2_1 _08515_ (.A(_02926_),
    .B(_02921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02927_));
 sky130_fd_sc_hd__a31o_1 _08516_ (.A1(_02916_),
    .A2(_02924_),
    .A3(_02925_),
    .B1(_02927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[4] ));
 sky130_fd_sc_hd__clkbuf_2 _08517_ (.A(_02898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02928_));
 sky130_fd_sc_hd__mux4_1 _08518_ (.A0(_02842_),
    .A1(_02858_),
    .A2(_02859_),
    .A3(_02860_),
    .S0(_02862_),
    .S1(_02863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02929_));
 sky130_fd_sc_hd__a22o_1 _08519_ (.A1(_02909_),
    .A2(_02920_),
    .B1(_02929_),
    .B2(_02867_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02930_));
 sky130_fd_sc_hd__and3_1 _08520_ (.A(_02857_),
    .B(_02919_),
    .C(_02929_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02931_));
 sky130_fd_sc_hd__nand2_2 _08521_ (.A(_02909_),
    .B(_02931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02932_));
 sky130_fd_sc_hd__and2_1 _08522_ (.A(_02930_),
    .B(_02932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02933_));
 sky130_fd_sc_hd__clkbuf_2 _08523_ (.A(_02933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02934_));
 sky130_fd_sc_hd__nand2_1 _08524_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[5] ),
    .B(_02934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02935_));
 sky130_fd_sc_hd__clkinv_2 _08525_ (.A(_02935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02936_));
 sky130_fd_sc_hd__nor2_1 _08526_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[5] ),
    .B(_02934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02937_));
 sky130_fd_sc_hd__or2_1 _08527_ (.A(_02936_),
    .B(_02937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02938_));
 sky130_fd_sc_hd__and2_1 _08528_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[4] ),
    .B(_02921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02939_));
 sky130_fd_sc_hd__inv_2 _08529_ (.A(_02939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02940_));
 sky130_fd_sc_hd__and2_1 _08530_ (.A(_02940_),
    .B(_02924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02941_));
 sky130_fd_sc_hd__xnor2_1 _08531_ (.A(_02938_),
    .B(_02941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02942_));
 sky130_fd_sc_hd__and3_1 _08532_ (.A(_02897_),
    .B(_02930_),
    .C(_02932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02943_));
 sky130_fd_sc_hd__o21bai_1 _08533_ (.A1(_02928_),
    .A2(_02942_),
    .B1_N(_02943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[5] ));
 sky130_fd_sc_hd__mux4_1 _08534_ (.A0(_02842_),
    .A1(_02880_),
    .A2(_02881_),
    .A3(_02885_),
    .S0(_02882_),
    .S1(_02863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02944_));
 sky130_fd_sc_hd__and2_2 _08535_ (.A(_02857_),
    .B(_02944_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02945_));
 sky130_fd_sc_hd__xnor2_4 _08536_ (.A(_02932_),
    .B(_02945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02946_));
 sky130_fd_sc_hd__clkbuf_2 _08537_ (.A(_02946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02947_));
 sky130_fd_sc_hd__xnor2_1 _08538_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[6] ),
    .B(_02946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02948_));
 sky130_fd_sc_hd__a311o_1 _08539_ (.A1(_02940_),
    .A2(_02924_),
    .A3(_02935_),
    .B1(_02937_),
    .C1(_02948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02949_));
 sky130_fd_sc_hd__clkbuf_4 _08540_ (.A(_02897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02950_));
 sky130_fd_sc_hd__o211a_1 _08541_ (.A1(_02937_),
    .A2(_02941_),
    .B1(_02948_),
    .C1(_02935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02951_));
 sky130_fd_sc_hd__nor2_1 _08542_ (.A(_02950_),
    .B(_02951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02952_));
 sky130_fd_sc_hd__a22o_1 _08543_ (.A1(_02928_),
    .A2(_02947_),
    .B1(_02949_),
    .B2(_02952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[6] ));
 sky130_fd_sc_hd__buf_2 _08544_ (.A(_02863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02953_));
 sky130_fd_sc_hd__mux2_1 _08545_ (.A0(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._00_ ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .S(_02886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02954_));
 sky130_fd_sc_hd__nor2_2 _08546_ (.A(_02882_),
    .B(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._00_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02955_));
 sky130_fd_sc_hd__o21ba_1 _08547_ (.A1(_02884_),
    .A2(_02954_),
    .B1_N(_02955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02956_));
 sky130_fd_sc_hd__inv_2 _08548_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02957_));
 sky130_fd_sc_hd__mux4_1 _08549_ (.A0(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .A2(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .A3(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ),
    .S0(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .S1(_02886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02958_));
 sky130_fd_sc_hd__or2_1 _08550_ (.A(_02957_),
    .B(_02958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02959_));
 sky130_fd_sc_hd__o211a_1 _08551_ (.A1(_02953_),
    .A2(_02956_),
    .B1(_02959_),
    .C1(_02857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02960_));
 sky130_fd_sc_hd__and3_1 _08552_ (.A(_02931_),
    .B(_02945_),
    .C(_02960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02961_));
 sky130_fd_sc_hd__nand2_1 _08553_ (.A(_02904_),
    .B(_02961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02962_));
 sky130_fd_sc_hd__a31o_1 _08554_ (.A1(_02904_),
    .A2(_02931_),
    .A3(_02945_),
    .B1(_02960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02963_));
 sky130_fd_sc_hd__and2_1 _08555_ (.A(_02962_),
    .B(_02963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02964_));
 sky130_fd_sc_hd__nor2_1 _08556_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[7] ),
    .B(_02964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02965_));
 sky130_fd_sc_hd__and3_1 _08557_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[7] ),
    .B(_02962_),
    .C(_02963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02966_));
 sky130_fd_sc_hd__or2_1 _08558_ (.A(_02965_),
    .B(_02966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02967_));
 sky130_fd_sc_hd__and2_1 _08559_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[6] ),
    .B(_02947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02968_));
 sky130_fd_sc_hd__or2b_1 _08560_ (.A(_02968_),
    .B_N(_02949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02969_));
 sky130_fd_sc_hd__xnor2_1 _08561_ (.A(_02967_),
    .B(_02969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02970_));
 sky130_fd_sc_hd__mux2_1 _08562_ (.A0(_02964_),
    .A1(_02970_),
    .S(_02914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02971_));
 sky130_fd_sc_hd__clkbuf_1 _08563_ (.A(_02971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[7] ));
 sky130_fd_sc_hd__or2_1 _08564_ (.A(_02957_),
    .B(_02849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02972_));
 sky130_fd_sc_hd__o21a_1 _08565_ (.A1(_02953_),
    .A2(_02842_),
    .B1(_02856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02973_));
 sky130_fd_sc_hd__and2_1 _08566_ (.A(_02972_),
    .B(_02973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02974_));
 sky130_fd_sc_hd__nand3_1 _08567_ (.A(_02904_),
    .B(_02961_),
    .C(_02974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02975_));
 sky130_fd_sc_hd__a21o_1 _08568_ (.A1(_02909_),
    .A2(_02961_),
    .B1(_02974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02976_));
 sky130_fd_sc_hd__and2_1 _08569_ (.A(_02975_),
    .B(_02976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02977_));
 sky130_fd_sc_hd__clkbuf_2 _08570_ (.A(_02977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02978_));
 sky130_fd_sc_hd__xnor2_1 _08571_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[8] ),
    .B(_02978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02979_));
 sky130_fd_sc_hd__nor2_1 _08572_ (.A(_02968_),
    .B(_02966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02980_));
 sky130_fd_sc_hd__a21o_1 _08573_ (.A1(_02949_),
    .A2(_02980_),
    .B1(_02965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02981_));
 sky130_fd_sc_hd__or2_1 _08574_ (.A(_02979_),
    .B(_02981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02982_));
 sky130_fd_sc_hd__a21oi_1 _08575_ (.A1(_02979_),
    .A2(_02981_),
    .B1(_02950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02983_));
 sky130_fd_sc_hd__a22o_1 _08576_ (.A1(_02928_),
    .A2(_02978_),
    .B1(_02982_),
    .B2(_02983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[8] ));
 sky130_fd_sc_hd__nand2_1 _08577_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[8] ),
    .B(_02978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02984_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08578_ (.A(_02957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02985_));
 sky130_fd_sc_hd__mux2_1 _08579_ (.A0(_02858_),
    .A1(_02859_),
    .S(_02882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02986_));
 sky130_fd_sc_hd__o21a_1 _08580_ (.A1(_02985_),
    .A2(_02986_),
    .B1(_02973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02987_));
 sky130_fd_sc_hd__and2_1 _08581_ (.A(_02972_),
    .B(_02987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02988_));
 sky130_fd_sc_hd__nand3_1 _08582_ (.A(_02903_),
    .B(_02961_),
    .C(_02988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02989_));
 sky130_fd_sc_hd__clkbuf_2 _08583_ (.A(_02989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02990_));
 sky130_fd_sc_hd__a31o_1 _08584_ (.A1(_02904_),
    .A2(_02961_),
    .A3(_02974_),
    .B1(_02987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02991_));
 sky130_fd_sc_hd__and3_1 _08585_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[9] ),
    .B(_02990_),
    .C(_02991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02992_));
 sky130_fd_sc_hd__a21oi_1 _08586_ (.A1(_02990_),
    .A2(_02991_),
    .B1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02993_));
 sky130_fd_sc_hd__or2_1 _08587_ (.A(_02992_),
    .B(_02993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02994_));
 sky130_fd_sc_hd__a21o_1 _08588_ (.A1(_02984_),
    .A2(_02982_),
    .B1(_02994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02995_));
 sky130_fd_sc_hd__nand2_1 _08589_ (.A(_02877_),
    .B(_02995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02996_));
 sky130_fd_sc_hd__and3_1 _08590_ (.A(_02984_),
    .B(_02982_),
    .C(_02994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02997_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08591_ (.A(_02990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02998_));
 sky130_fd_sc_hd__and2_1 _08592_ (.A(_02998_),
    .B(_02991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02999_));
 sky130_fd_sc_hd__a2bb2o_1 _08593_ (.A1_N(_02996_),
    .A2_N(_02997_),
    .B1(_02999_),
    .B2(_02928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[9] ));
 sky130_fd_sc_hd__o21ai_2 _08594_ (.A1(_02953_),
    .A2(_02843_),
    .B1(_02867_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03000_));
 sky130_fd_sc_hd__nor2_1 _08595_ (.A(_02985_),
    .B(_02883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03001_));
 sky130_fd_sc_hd__nor2_1 _08596_ (.A(_03000_),
    .B(_03001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03002_));
 sky130_fd_sc_hd__xnor2_1 _08597_ (.A(_02989_),
    .B(_03002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03003_));
 sky130_fd_sc_hd__xnor2_1 _08598_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[10] ),
    .B(_03003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03004_));
 sky130_fd_sc_hd__a21oi_1 _08599_ (.A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[8] ),
    .A2(_02978_),
    .B1(_02992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03005_));
 sky130_fd_sc_hd__a21o_1 _08600_ (.A1(_02982_),
    .A2(_03005_),
    .B1(_02993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03006_));
 sky130_fd_sc_hd__xor2_1 _08601_ (.A(_03004_),
    .B(_03006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03007_));
 sky130_fd_sc_hd__clkbuf_2 _08602_ (.A(_03003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03008_));
 sky130_fd_sc_hd__and2_1 _08603_ (.A(_02898_),
    .B(_03008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03009_));
 sky130_fd_sc_hd__a21o_1 _08604_ (.A1(_02878_),
    .A2(_03007_),
    .B1(_03009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[10] ));
 sky130_fd_sc_hd__inv_2 _08605_ (.A(_03002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03010_));
 sky130_fd_sc_hd__nor2_2 _08606_ (.A(_02985_),
    .B(_02900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03011_));
 sky130_fd_sc_hd__or3_1 _08607_ (.A(_02989_),
    .B(_03010_),
    .C(_03011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03012_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08608_ (.A(_03012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03013_));
 sky130_fd_sc_hd__o22ai_4 _08609_ (.A1(_02990_),
    .A2(_03010_),
    .B1(_03011_),
    .B2(_03000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03014_));
 sky130_fd_sc_hd__and3_1 _08610_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[11] ),
    .B(_03013_),
    .C(_03014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03015_));
 sky130_fd_sc_hd__a21oi_1 _08611_ (.A1(_03013_),
    .A2(_03014_),
    .B1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03016_));
 sky130_fd_sc_hd__or2_1 _08612_ (.A(_03015_),
    .B(_03016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03017_));
 sky130_fd_sc_hd__o2bb2ai_1 _08613_ (.A1_N(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[10] ),
    .A2_N(_03008_),
    .B1(_03004_),
    .B2(_03006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03018_));
 sky130_fd_sc_hd__xnor2_1 _08614_ (.A(_03017_),
    .B(_03018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03019_));
 sky130_fd_sc_hd__and3_1 _08615_ (.A(_02926_),
    .B(_03013_),
    .C(_03014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03020_));
 sky130_fd_sc_hd__a21o_1 _08616_ (.A1(_02878_),
    .A2(_03019_),
    .B1(_03020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[11] ));
 sky130_fd_sc_hd__clkbuf_2 _08617_ (.A(_02854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03021_));
 sky130_fd_sc_hd__a21o_1 _08618_ (.A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[10] ),
    .A2(_03008_),
    .B1(_03015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03022_));
 sky130_fd_sc_hd__or2b_1 _08619_ (.A(_03016_),
    .B_N(_03022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03023_));
 sky130_fd_sc_hd__or3_1 _08620_ (.A(_03004_),
    .B(_03015_),
    .C(_03016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03024_));
 sky130_fd_sc_hd__or3_1 _08621_ (.A(_02993_),
    .B(_03005_),
    .C(_03024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03025_));
 sky130_fd_sc_hd__or2_1 _08622_ (.A(_02979_),
    .B(_02994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03026_));
 sky130_fd_sc_hd__a2111o_1 _08623_ (.A1(_02949_),
    .A2(_02980_),
    .B1(_03024_),
    .C1(_03026_),
    .D1(_02965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03027_));
 sky130_fd_sc_hd__o21ba_1 _08624_ (.A1(_02884_),
    .A2(_02917_),
    .B1_N(_02955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03028_));
 sky130_fd_sc_hd__o31a_1 _08625_ (.A1(_02998_),
    .A2(_03001_),
    .A3(_03011_),
    .B1(_02973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03029_));
 sky130_fd_sc_hd__o21a_1 _08626_ (.A1(_02985_),
    .A2(_03028_),
    .B1(_03029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03030_));
 sky130_fd_sc_hd__clkbuf_2 _08627_ (.A(_03030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03031_));
 sky130_fd_sc_hd__xnor2_1 _08628_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[12] ),
    .B(_03031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03032_));
 sky130_fd_sc_hd__a31o_1 _08629_ (.A1(_03023_),
    .A2(_03025_),
    .A3(_03027_),
    .B1(_03032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03033_));
 sky130_fd_sc_hd__nand4_1 _08630_ (.A(_03032_),
    .B(_03023_),
    .C(_03025_),
    .D(_03027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03034_));
 sky130_fd_sc_hd__and2_1 _08631_ (.A(_02926_),
    .B(_03031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03035_));
 sky130_fd_sc_hd__a31o_1 _08632_ (.A1(_03021_),
    .A2(_03033_),
    .A3(_03034_),
    .B1(_03035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[12] ));
 sky130_fd_sc_hd__clkbuf_2 _08633_ (.A(_02877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03036_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08634_ (.A(_03029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03037_));
 sky130_fd_sc_hd__nor2_1 _08635_ (.A(_02884_),
    .B(_02858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03038_));
 sky130_fd_sc_hd__o21ai_4 _08636_ (.A1(_02955_),
    .A2(_03038_),
    .B1(_02953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03039_));
 sky130_fd_sc_hd__and3_1 _08637_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[13] ),
    .B(_03037_),
    .C(_03039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03040_));
 sky130_fd_sc_hd__a21oi_1 _08638_ (.A1(_03037_),
    .A2(_03039_),
    .B1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03041_));
 sky130_fd_sc_hd__or2_1 _08639_ (.A(_03040_),
    .B(_03041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03042_));
 sky130_fd_sc_hd__a21bo_1 _08640_ (.A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[12] ),
    .A2(_03031_),
    .B1_N(_03033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03043_));
 sky130_fd_sc_hd__xnor2_1 _08641_ (.A(_03042_),
    .B(_03043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03044_));
 sky130_fd_sc_hd__and3_1 _08642_ (.A(_02898_),
    .B(_03037_),
    .C(_03039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03045_));
 sky130_fd_sc_hd__a21o_1 _08643_ (.A1(_03036_),
    .A2(_03044_),
    .B1(_03045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[13] ));
 sky130_fd_sc_hd__nor2_1 _08644_ (.A(_03040_),
    .B(_03043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03046_));
 sky130_fd_sc_hd__nor2_1 _08645_ (.A(_02884_),
    .B(_02880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03047_));
 sky130_fd_sc_hd__o21ai_1 _08646_ (.A1(_02955_),
    .A2(_03047_),
    .B1(_02953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03048_));
 sky130_fd_sc_hd__o311a_1 _08647_ (.A1(_02990_),
    .A2(_03001_),
    .A3(_03011_),
    .B1(_03048_),
    .C1(_02973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03049_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08648_ (.A(_03049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03050_));
 sky130_fd_sc_hd__nand2_1 _08649_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[14] ),
    .B(_03050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03051_));
 sky130_fd_sc_hd__or2_1 _08650_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[14] ),
    .B(_03049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03052_));
 sky130_fd_sc_hd__nand2_1 _08651_ (.A(_03051_),
    .B(_03052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03053_));
 sky130_fd_sc_hd__o21ai_1 _08652_ (.A1(_03041_),
    .A2(_03046_),
    .B1(_03053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03054_));
 sky130_fd_sc_hd__or2_1 _08653_ (.A(_03041_),
    .B(_03053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03055_));
 sky130_fd_sc_hd__or2_1 _08654_ (.A(_03046_),
    .B(_03055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03056_));
 sky130_fd_sc_hd__and2_1 _08655_ (.A(_02926_),
    .B(_03050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03057_));
 sky130_fd_sc_hd__a31o_1 _08656_ (.A1(_03021_),
    .A2(_03054_),
    .A3(_03056_),
    .B1(_03057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[14] ));
 sky130_fd_sc_hd__or2_1 _08657_ (.A(_02985_),
    .B(_02956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03058_));
 sky130_fd_sc_hd__o311a_2 _08658_ (.A1(_02998_),
    .A2(_03001_),
    .A3(_03011_),
    .B1(_03058_),
    .C1(_02973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03059_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08659_ (.A(_03059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03060_));
 sky130_fd_sc_hd__and2_1 _08660_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[15] ),
    .B(_03060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03061_));
 sky130_fd_sc_hd__nor2_1 _08661_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[15] ),
    .B(_03060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03062_));
 sky130_fd_sc_hd__or2_2 _08662_ (.A(_03061_),
    .B(_03062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03063_));
 sky130_fd_sc_hd__a21o_1 _08663_ (.A1(_03051_),
    .A2(_03056_),
    .B1(_03063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03064_));
 sky130_fd_sc_hd__nand3_1 _08664_ (.A(_03051_),
    .B(_03056_),
    .C(_03063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03065_));
 sky130_fd_sc_hd__and2_1 _08665_ (.A(_02926_),
    .B(_03060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03066_));
 sky130_fd_sc_hd__a31o_1 _08666_ (.A1(_03021_),
    .A2(_03064_),
    .A3(_03065_),
    .B1(_03066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[15] ));
 sky130_fd_sc_hd__a21oi_1 _08667_ (.A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[12] ),
    .A2(_03031_),
    .B1(_03040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03067_));
 sky130_fd_sc_hd__a21oi_1 _08668_ (.A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[14] ),
    .A2(_03050_),
    .B1(_03061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03068_));
 sky130_fd_sc_hd__o32a_1 _08669_ (.A1(_03067_),
    .A2(_03055_),
    .A3(_03063_),
    .B1(_03068_),
    .B2(_03062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03069_));
 sky130_fd_sc_hd__o41ai_4 _08670_ (.A1(_03033_),
    .A2(_03042_),
    .A3(_03053_),
    .A4(_03063_),
    .B1(_03069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03070_));
 sky130_fd_sc_hd__and3_2 _08671_ (.A(_02867_),
    .B(_02843_),
    .C(_03012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03071_));
 sky130_fd_sc_hd__clkbuf_2 _08672_ (.A(_03071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03072_));
 sky130_fd_sc_hd__clkbuf_2 _08673_ (.A(_03072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03073_));
 sky130_fd_sc_hd__xnor2_1 _08674_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[16] ),
    .B(_03073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03074_));
 sky130_fd_sc_hd__xnor2_1 _08675_ (.A(_03070_),
    .B(_03074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03075_));
 sky130_fd_sc_hd__clkbuf_2 _08676_ (.A(_03071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03076_));
 sky130_fd_sc_hd__clkbuf_2 _08677_ (.A(_03076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03077_));
 sky130_fd_sc_hd__buf_2 _08678_ (.A(_03077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03078_));
 sky130_fd_sc_hd__buf_2 _08679_ (.A(_03078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03079_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08680_ (.A(_03079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03080_));
 sky130_fd_sc_hd__clkbuf_2 _08681_ (.A(_03080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03081_));
 sky130_fd_sc_hd__and2_1 _08682_ (.A(_02896_),
    .B(_03081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03082_));
 sky130_fd_sc_hd__clkbuf_2 _08683_ (.A(_03082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03083_));
 sky130_fd_sc_hd__clkbuf_2 _08684_ (.A(_03083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03084_));
 sky130_fd_sc_hd__a21o_1 _08685_ (.A1(_03036_),
    .A2(_03075_),
    .B1(_03084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[16] ));
 sky130_fd_sc_hd__clkbuf_2 _08686_ (.A(_03078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03085_));
 sky130_fd_sc_hd__clkbuf_2 _08687_ (.A(_03085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03086_));
 sky130_fd_sc_hd__clkbuf_2 _08688_ (.A(_03086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03087_));
 sky130_fd_sc_hd__and2b_1 _08689_ (.A_N(_03074_),
    .B(_03070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03088_));
 sky130_fd_sc_hd__a21oi_1 _08690_ (.A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[16] ),
    .A2(_03087_),
    .B1(_03088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03089_));
 sky130_fd_sc_hd__nand2_1 _08691_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[17] ),
    .B(_03073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03090_));
 sky130_fd_sc_hd__or2_1 _08692_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[17] ),
    .B(_03076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03091_));
 sky130_fd_sc_hd__nand2_1 _08693_ (.A(_03090_),
    .B(_03091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03092_));
 sky130_fd_sc_hd__or2_1 _08694_ (.A(_03089_),
    .B(_03092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03093_));
 sky130_fd_sc_hd__nand2_1 _08695_ (.A(_03089_),
    .B(_03092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03094_));
 sky130_fd_sc_hd__clkbuf_2 _08696_ (.A(_03083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03095_));
 sky130_fd_sc_hd__a31o_1 _08697_ (.A1(_03021_),
    .A2(_03093_),
    .A3(_03094_),
    .B1(_03095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[17] ));
 sky130_fd_sc_hd__or2b_1 _08698_ (.A(_03089_),
    .B_N(_03091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03096_));
 sky130_fd_sc_hd__nand2_1 _08699_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[18] ),
    .B(_03073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03097_));
 sky130_fd_sc_hd__clkbuf_2 _08700_ (.A(_03071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03098_));
 sky130_fd_sc_hd__or2_1 _08701_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[18] ),
    .B(_03098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03099_));
 sky130_fd_sc_hd__nand2_1 _08702_ (.A(_03097_),
    .B(_03099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03100_));
 sky130_fd_sc_hd__a21o_1 _08703_ (.A1(_03090_),
    .A2(_03096_),
    .B1(_03100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03101_));
 sky130_fd_sc_hd__nand3_1 _08704_ (.A(_03090_),
    .B(_03096_),
    .C(_03100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03102_));
 sky130_fd_sc_hd__a31o_1 _08705_ (.A1(_03021_),
    .A2(_03101_),
    .A3(_03102_),
    .B1(_03095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[18] ));
 sky130_fd_sc_hd__clkbuf_2 _08706_ (.A(_02875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03103_));
 sky130_fd_sc_hd__xnor2_1 _08707_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[19] ),
    .B(_03073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03104_));
 sky130_fd_sc_hd__a21o_1 _08708_ (.A1(_03097_),
    .A2(_03101_),
    .B1(_03104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03105_));
 sky130_fd_sc_hd__nand3_1 _08709_ (.A(_03097_),
    .B(_03101_),
    .C(_03104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03106_));
 sky130_fd_sc_hd__a31o_1 _08710_ (.A1(_03103_),
    .A2(_03105_),
    .A3(_03106_),
    .B1(_03095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[19] ));
 sky130_fd_sc_hd__nand2_1 _08711_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[20] ),
    .B(_03077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03107_));
 sky130_fd_sc_hd__or2_1 _08712_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[20] ),
    .B(_03098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03108_));
 sky130_fd_sc_hd__nand2_1 _08713_ (.A(_03107_),
    .B(_03108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03109_));
 sky130_fd_sc_hd__or4_1 _08714_ (.A(_03074_),
    .B(_03092_),
    .C(_03100_),
    .D(_03104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03110_));
 sky130_fd_sc_hd__inv_2 _08715_ (.A(_03110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03111_));
 sky130_fd_sc_hd__o41a_1 _08716_ (.A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[16] ),
    .A2(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[17] ),
    .A3(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[18] ),
    .A4(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[19] ),
    .B1(_03078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03112_));
 sky130_fd_sc_hd__a21oi_1 _08717_ (.A1(_03070_),
    .A2(_03111_),
    .B1(_03112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03113_));
 sky130_fd_sc_hd__xor2_1 _08718_ (.A(_03109_),
    .B(_03113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03114_));
 sky130_fd_sc_hd__a21o_1 _08719_ (.A1(_03036_),
    .A2(_03114_),
    .B1(_03084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[20] ));
 sky130_fd_sc_hd__o21a_1 _08720_ (.A1(_03109_),
    .A2(_03113_),
    .B1(_03107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03115_));
 sky130_fd_sc_hd__nand2_1 _08721_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[21] ),
    .B(_03077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03116_));
 sky130_fd_sc_hd__buf_2 _08722_ (.A(_03071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03117_));
 sky130_fd_sc_hd__or2_1 _08723_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[21] ),
    .B(_03117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03118_));
 sky130_fd_sc_hd__nand2_1 _08724_ (.A(_03116_),
    .B(_03118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03119_));
 sky130_fd_sc_hd__or2_1 _08725_ (.A(_03115_),
    .B(_03119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03120_));
 sky130_fd_sc_hd__nand2_1 _08726_ (.A(_03115_),
    .B(_03119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03121_));
 sky130_fd_sc_hd__a31o_1 _08727_ (.A1(_03103_),
    .A2(_03120_),
    .A3(_03121_),
    .B1(_03095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[21] ));
 sky130_fd_sc_hd__or2b_1 _08728_ (.A(_03115_),
    .B_N(_03118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03122_));
 sky130_fd_sc_hd__and2_1 _08729_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[22] ),
    .B(_03076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03123_));
 sky130_fd_sc_hd__nor2_1 _08730_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[22] ),
    .B(_03073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03124_));
 sky130_fd_sc_hd__or2_1 _08731_ (.A(_03123_),
    .B(_03124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03125_));
 sky130_fd_sc_hd__a21oi_1 _08732_ (.A1(_03116_),
    .A2(_03122_),
    .B1(_03125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03126_));
 sky130_fd_sc_hd__clkbuf_2 _08733_ (.A(_02897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03127_));
 sky130_fd_sc_hd__a31o_1 _08734_ (.A1(_03116_),
    .A2(_03122_),
    .A3(_03125_),
    .B1(_03127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03128_));
 sky130_fd_sc_hd__clkbuf_2 _08735_ (.A(_03082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03129_));
 sky130_fd_sc_hd__o21bai_1 _08736_ (.A1(_03126_),
    .A2(_03128_),
    .B1_N(_03129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[22] ));
 sky130_fd_sc_hd__xor2_1 _08737_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[23] ),
    .B(_03077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03130_));
 sky130_fd_sc_hd__o21ai_1 _08738_ (.A1(_03123_),
    .A2(_03126_),
    .B1(_03130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03131_));
 sky130_fd_sc_hd__or3_1 _08739_ (.A(_03123_),
    .B(_03126_),
    .C(_03130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03132_));
 sky130_fd_sc_hd__a31o_1 _08740_ (.A1(_03103_),
    .A2(_03131_),
    .A3(_03132_),
    .B1(_03095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[23] ));
 sky130_fd_sc_hd__or4b_1 _08741_ (.A(_03109_),
    .B(_03119_),
    .C(_03125_),
    .D_N(_03130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03133_));
 sky130_fd_sc_hd__nor2_1 _08742_ (.A(_03110_),
    .B(_03133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03134_));
 sky130_fd_sc_hd__o41a_1 _08743_ (.A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[20] ),
    .A2(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[21] ),
    .A3(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[22] ),
    .A4(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[23] ),
    .B1(_03078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03135_));
 sky130_fd_sc_hd__or2_1 _08744_ (.A(_03112_),
    .B(_03135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03136_));
 sky130_fd_sc_hd__a21o_1 _08745_ (.A1(_03070_),
    .A2(_03134_),
    .B1(_03136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03137_));
 sky130_fd_sc_hd__buf_2 _08746_ (.A(_03077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03138_));
 sky130_fd_sc_hd__xor2_1 _08747_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[24] ),
    .B(_03138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03139_));
 sky130_fd_sc_hd__nand2_1 _08748_ (.A(_03137_),
    .B(_03139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03140_));
 sky130_fd_sc_hd__o21a_1 _08749_ (.A1(_03137_),
    .A2(_03139_),
    .B1(_02877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03141_));
 sky130_fd_sc_hd__a21o_1 _08750_ (.A1(_03140_),
    .A2(_03141_),
    .B1(_03084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[24] ));
 sky130_fd_sc_hd__xor2_1 _08751_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[25] ),
    .B(_03138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03142_));
 sky130_fd_sc_hd__buf_2 _08752_ (.A(_03087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03143_));
 sky130_fd_sc_hd__a22o_1 _08753_ (.A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[24] ),
    .A2(_03143_),
    .B1(_03137_),
    .B2(_03139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03144_));
 sky130_fd_sc_hd__xor2_1 _08754_ (.A(_03142_),
    .B(_03144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03145_));
 sky130_fd_sc_hd__a21o_1 _08755_ (.A1(_03036_),
    .A2(_03145_),
    .B1(_03084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[25] ));
 sky130_fd_sc_hd__o21ai_1 _08756_ (.A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[24] ),
    .A2(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[25] ),
    .B1(_03081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03146_));
 sky130_fd_sc_hd__and2_1 _08757_ (.A(_03139_),
    .B(_03142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03147_));
 sky130_fd_sc_hd__nand2_1 _08758_ (.A(_03137_),
    .B(_03147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03148_));
 sky130_fd_sc_hd__nand2_1 _08759_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[26] ),
    .B(_03085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03149_));
 sky130_fd_sc_hd__or2_1 _08760_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[26] ),
    .B(_03138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03150_));
 sky130_fd_sc_hd__nand2_1 _08761_ (.A(_03149_),
    .B(_03150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03151_));
 sky130_fd_sc_hd__a21o_1 _08762_ (.A1(_03146_),
    .A2(_03148_),
    .B1(_03151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03152_));
 sky130_fd_sc_hd__nand3_1 _08763_ (.A(_03151_),
    .B(_03146_),
    .C(_03148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03153_));
 sky130_fd_sc_hd__buf_2 _08764_ (.A(_03082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03154_));
 sky130_fd_sc_hd__a31o_1 _08765_ (.A1(_03103_),
    .A2(_03152_),
    .A3(_03153_),
    .B1(_03154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[26] ));
 sky130_fd_sc_hd__xnor2_1 _08766_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[27] ),
    .B(_03085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03155_));
 sky130_fd_sc_hd__nand2_1 _08767_ (.A(_03149_),
    .B(_03152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03156_));
 sky130_fd_sc_hd__xnor2_1 _08768_ (.A(_03155_),
    .B(_03156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03157_));
 sky130_fd_sc_hd__a21o_1 _08769_ (.A1(_03036_),
    .A2(_03157_),
    .B1(_03084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[27] ));
 sky130_fd_sc_hd__nor2_1 _08770_ (.A(_03151_),
    .B(_03155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03158_));
 sky130_fd_sc_hd__o41a_1 _08771_ (.A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[24] ),
    .A2(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[25] ),
    .A3(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[26] ),
    .A4(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[27] ),
    .B1(_03086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03159_));
 sky130_fd_sc_hd__a31oi_2 _08772_ (.A1(_03137_),
    .A2(_03147_),
    .A3(_03158_),
    .B1(_03159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03160_));
 sky130_fd_sc_hd__and2_1 _08773_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[28] ),
    .B(_03079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03161_));
 sky130_fd_sc_hd__nor2_1 _08774_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[28] ),
    .B(_03086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03162_));
 sky130_fd_sc_hd__or2_1 _08775_ (.A(_03161_),
    .B(_03162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03163_));
 sky130_fd_sc_hd__nor2_1 _08776_ (.A(_03160_),
    .B(_03163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03164_));
 sky130_fd_sc_hd__a21o_1 _08777_ (.A1(_03160_),
    .A2(_03163_),
    .B1(_02950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03165_));
 sky130_fd_sc_hd__o21bai_1 _08778_ (.A1(_03164_),
    .A2(_03165_),
    .B1_N(_03129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[28] ));
 sky130_fd_sc_hd__nand2_1 _08779_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[29] ),
    .B(_03080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03166_));
 sky130_fd_sc_hd__or2_1 _08780_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[29] ),
    .B(_03080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03167_));
 sky130_fd_sc_hd__o211ai_1 _08781_ (.A1(_03161_),
    .A2(_03164_),
    .B1(_03166_),
    .C1(_03167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03168_));
 sky130_fd_sc_hd__a211o_1 _08782_ (.A1(_03166_),
    .A2(_03167_),
    .B1(_03161_),
    .C1(_03164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03169_));
 sky130_fd_sc_hd__a31o_1 _08783_ (.A1(_03103_),
    .A2(_03168_),
    .A3(_03169_),
    .B1(_03154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[29] ));
 sky130_fd_sc_hd__buf_2 _08784_ (.A(_02875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03170_));
 sky130_fd_sc_hd__o21ai_1 _08785_ (.A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[28] ),
    .A2(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[29] ),
    .B1(_03143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03171_));
 sky130_fd_sc_hd__or4bb_1 _08786_ (.A(_03160_),
    .B(_03163_),
    .C_N(_03166_),
    .D_N(_03167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03172_));
 sky130_fd_sc_hd__nand2_1 _08787_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[30] ),
    .B(_03081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03173_));
 sky130_fd_sc_hd__or2_1 _08788_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[30] ),
    .B(_03087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03174_));
 sky130_fd_sc_hd__nand2_1 _08789_ (.A(_03173_),
    .B(_03174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03175_));
 sky130_fd_sc_hd__a21o_1 _08790_ (.A1(_03171_),
    .A2(_03172_),
    .B1(_03175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03176_));
 sky130_fd_sc_hd__nand3_1 _08791_ (.A(_03175_),
    .B(_03171_),
    .C(_03172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03177_));
 sky130_fd_sc_hd__a31o_1 _08792_ (.A1(_03170_),
    .A2(_03176_),
    .A3(_03177_),
    .B1(_03154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[30] ));
 sky130_fd_sc_hd__xnor2_1 _08793_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[31] ),
    .B(_03143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03178_));
 sky130_fd_sc_hd__a21oi_1 _08794_ (.A1(_03173_),
    .A2(_03176_),
    .B1(_03178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03179_));
 sky130_fd_sc_hd__a31o_1 _08795_ (.A1(_03173_),
    .A2(_03176_),
    .A3(_03178_),
    .B1(_03127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03180_));
 sky130_fd_sc_hd__o21bai_1 _08796_ (.A1(_03179_),
    .A2(_03180_),
    .B1_N(_03129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[31] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08797_ (.A(\sa_inst.sak._13_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03181_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08798_ (.A(_03181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03182_));
 sky130_fd_sc_hd__clkbuf_1 _08799_ (.A(\sa_inst.sak._03_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03183_));
 sky130_fd_sc_hd__nand2_1 _08800_ (.A(_03182_),
    .B(_03183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03184_));
 sky130_fd_sc_hd__xnor2_1 _08801_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._01_ ),
    .B(_03184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03185_));
 sky130_fd_sc_hd__clkbuf_2 _08802_ (.A(\sa_inst.sak._03_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03186_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08803_ (.A(\sa_inst.sak._13_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03187_));
 sky130_fd_sc_hd__a22oi_1 _08804_ (.A1(_03182_),
    .A2(_03186_),
    .B1(_03187_),
    .B2(_03183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03188_));
 sky130_fd_sc_hd__and2_1 _08805_ (.A(\sa_inst.sak._03_[5] ),
    .B(_03187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03189_));
 sky130_fd_sc_hd__and3_1 _08806_ (.A(_03182_),
    .B(_03183_),
    .C(_03189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03190_));
 sky130_fd_sc_hd__or2_1 _08807_ (.A(_03188_),
    .B(_03190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03191_));
 sky130_fd_sc_hd__xnor2_1 _08808_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._01_ ),
    .B(_03191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03192_));
 sky130_fd_sc_hd__xor2_4 _08809_ (.A(_02672_),
    .B(\sa_inst.sak._03_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03193_));
 sky130_fd_sc_hd__clkbuf_2 _08810_ (.A(_03193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03194_));
 sky130_fd_sc_hd__mux2_1 _08811_ (.A0(_03185_),
    .A1(_03192_),
    .S(_03194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03195_));
 sky130_fd_sc_hd__clkbuf_1 _08812_ (.A(_03195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[1] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08813_ (.A(\sa_inst.sak._03_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03196_));
 sky130_fd_sc_hd__and3_1 _08814_ (.A(_03181_),
    .B(_03196_),
    .C(_03189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03197_));
 sky130_fd_sc_hd__a21oi_1 _08815_ (.A1(_03182_),
    .A2(_03196_),
    .B1(_03189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03198_));
 sky130_fd_sc_hd__nor2_1 _08816_ (.A(_03197_),
    .B(_03198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03199_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08817_ (.A(\sa_inst.sak._13_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03200_));
 sky130_fd_sc_hd__clkbuf_2 _08818_ (.A(_03200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03201_));
 sky130_fd_sc_hd__nand2_1 _08819_ (.A(_03183_),
    .B(_03201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03202_));
 sky130_fd_sc_hd__xnor2_1 _08820_ (.A(_03199_),
    .B(_03202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03203_));
 sky130_fd_sc_hd__xnor2_1 _08821_ (.A(_03190_),
    .B(_03203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03204_));
 sky130_fd_sc_hd__xnor2_1 _08822_ (.A(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._01_ ),
    .B(_03204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03205_));
 sky130_fd_sc_hd__mux2_1 _08823_ (.A0(_03192_),
    .A1(_03205_),
    .S(_03194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03206_));
 sky130_fd_sc_hd__clkbuf_1 _08824_ (.A(_03206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[2] ));
 sky130_fd_sc_hd__buf_2 _08825_ (.A(_02841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03207_));
 sky130_fd_sc_hd__and2_1 _08826_ (.A(_03190_),
    .B(_03203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03208_));
 sky130_fd_sc_hd__clkbuf_2 _08827_ (.A(\sa_inst.sak._03_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03209_));
 sky130_fd_sc_hd__nand2_1 _08828_ (.A(_03182_),
    .B(_03209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03210_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08829_ (.A(\sa_inst.sak._13_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03211_));
 sky130_fd_sc_hd__clkbuf_2 _08830_ (.A(_03211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03212_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08831_ (.A(\sa_inst.sak._03_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03213_));
 sky130_fd_sc_hd__a22oi_1 _08832_ (.A1(_03187_),
    .A2(_03213_),
    .B1(_03201_),
    .B2(_03186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03214_));
 sky130_fd_sc_hd__and3_1 _08833_ (.A(_03213_),
    .B(_03201_),
    .C(_03189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03215_));
 sky130_fd_sc_hd__o2bb2a_1 _08834_ (.A1_N(_03183_),
    .A2_N(_03212_),
    .B1(_03214_),
    .B2(_03215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03216_));
 sky130_fd_sc_hd__and4bb_1 _08835_ (.A_N(_03214_),
    .B_N(_03215_),
    .C(\sa_inst.sak._03_[4] ),
    .D(_03212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03217_));
 sky130_fd_sc_hd__nor2_1 _08836_ (.A(_03216_),
    .B(_03217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03218_));
 sky130_fd_sc_hd__xnor2_1 _08837_ (.A(_03210_),
    .B(_03218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03219_));
 sky130_fd_sc_hd__o21ba_1 _08838_ (.A1(_03198_),
    .A2(_03202_),
    .B1_N(_03197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03220_));
 sky130_fd_sc_hd__xnor2_1 _08839_ (.A(_03219_),
    .B(_03220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03221_));
 sky130_fd_sc_hd__and2_1 _08840_ (.A(_03208_),
    .B(_03221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03222_));
 sky130_fd_sc_hd__nor2_1 _08841_ (.A(_03208_),
    .B(_03221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03223_));
 sky130_fd_sc_hd__or2_1 _08842_ (.A(_03222_),
    .B(_03223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03224_));
 sky130_fd_sc_hd__xnor2_1 _08843_ (.A(_03207_),
    .B(_03224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03225_));
 sky130_fd_sc_hd__mux2_1 _08844_ (.A0(_03205_),
    .A1(_03225_),
    .S(_03194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03226_));
 sky130_fd_sc_hd__clkbuf_1 _08845_ (.A(_03226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[3] ));
 sky130_fd_sc_hd__and2b_1 _08846_ (.A_N(_03220_),
    .B(_03219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03227_));
 sky130_fd_sc_hd__or3_1 _08847_ (.A(_03210_),
    .B(_03216_),
    .C(_03217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03228_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08848_ (.A(\sa_inst.sak._03_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03229_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08849_ (.A(_03229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03230_));
 sky130_fd_sc_hd__a22oi_1 _08850_ (.A1(_03187_),
    .A2(_03209_),
    .B1(_03230_),
    .B2(_03181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03231_));
 sky130_fd_sc_hd__and4_1 _08851_ (.A(_03181_),
    .B(_03187_),
    .C(\sa_inst.sak._03_[7] ),
    .D(_03229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03232_));
 sky130_fd_sc_hd__nor2_1 _08852_ (.A(_03231_),
    .B(_03232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03233_));
 sky130_fd_sc_hd__a22oi_1 _08853_ (.A1(_03213_),
    .A2(_03200_),
    .B1(_03211_),
    .B2(\sa_inst.sak._03_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03234_));
 sky130_fd_sc_hd__and4_1 _08854_ (.A(\sa_inst.sak._03_[5] ),
    .B(\sa_inst.sak._03_[6] ),
    .C(_03200_),
    .D(\sa_inst.sak._13_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03235_));
 sky130_fd_sc_hd__nor2_1 _08855_ (.A(_03234_),
    .B(_03235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03236_));
 sky130_fd_sc_hd__nand2_1 _08856_ (.A(\sa_inst.sak._03_[4] ),
    .B(\sa_inst.sak._13_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03237_));
 sky130_fd_sc_hd__xnor2_1 _08857_ (.A(_03236_),
    .B(_03237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03238_));
 sky130_fd_sc_hd__xnor2_1 _08858_ (.A(_03233_),
    .B(_03238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03239_));
 sky130_fd_sc_hd__and2_1 _08859_ (.A(_03228_),
    .B(_03239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03240_));
 sky130_fd_sc_hd__nor2_1 _08860_ (.A(_03228_),
    .B(_03239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03241_));
 sky130_fd_sc_hd__nor2_1 _08861_ (.A(_03240_),
    .B(_03241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03242_));
 sky130_fd_sc_hd__or2_1 _08862_ (.A(_03215_),
    .B(_03217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03243_));
 sky130_fd_sc_hd__xor2_1 _08863_ (.A(_03242_),
    .B(_03243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03244_));
 sky130_fd_sc_hd__o21ai_2 _08864_ (.A1(_03227_),
    .A2(_03222_),
    .B1(_03244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03245_));
 sky130_fd_sc_hd__or3_1 _08865_ (.A(_03227_),
    .B(_03222_),
    .C(_03244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03246_));
 sky130_fd_sc_hd__nand2_1 _08866_ (.A(_03245_),
    .B(_03246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03247_));
 sky130_fd_sc_hd__xnor2_1 _08867_ (.A(_03207_),
    .B(_03247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03248_));
 sky130_fd_sc_hd__mux2_1 _08868_ (.A0(_03225_),
    .A1(_03248_),
    .S(_03194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03249_));
 sky130_fd_sc_hd__clkbuf_1 _08869_ (.A(_03249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[4] ));
 sky130_fd_sc_hd__and2_1 _08870_ (.A(_03233_),
    .B(_03238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03250_));
 sky130_fd_sc_hd__a22oi_1 _08871_ (.A1(\sa_inst.sak._13_[5] ),
    .A2(\sa_inst.sak._03_[8] ),
    .B1(\sa_inst.sak._03_[9] ),
    .B2(_03181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03251_));
 sky130_fd_sc_hd__and4_1 _08872_ (.A(\sa_inst.sak._13_[4] ),
    .B(\sa_inst.sak._13_[5] ),
    .C(\sa_inst.sak._03_[8] ),
    .D(\sa_inst.sak._03_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03252_));
 sky130_fd_sc_hd__o2bb2a_1 _08873_ (.A1_N(_03200_),
    .A2_N(\sa_inst.sak._03_[7] ),
    .B1(_03251_),
    .B2(_03252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03253_));
 sky130_fd_sc_hd__and4bb_1 _08874_ (.A_N(_03251_),
    .B_N(_03252_),
    .C(_03200_),
    .D(\sa_inst.sak._03_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03254_));
 sky130_fd_sc_hd__nor2_1 _08875_ (.A(_03253_),
    .B(_03254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03255_));
 sky130_fd_sc_hd__xnor2_1 _08876_ (.A(_03232_),
    .B(_03255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03256_));
 sky130_fd_sc_hd__a22oi_2 _08877_ (.A1(_03213_),
    .A2(_03211_),
    .B1(\sa_inst.sak._13_[8] ),
    .B2(_03186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03257_));
 sky130_fd_sc_hd__and4_2 _08878_ (.A(\sa_inst.sak._03_[5] ),
    .B(\sa_inst.sak._03_[6] ),
    .C(_03211_),
    .D(\sa_inst.sak._13_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03258_));
 sky130_fd_sc_hd__nand2_1 _08879_ (.A(\sa_inst.sak._03_[4] ),
    .B(\sa_inst.sak._13_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03259_));
 sky130_fd_sc_hd__o21a_1 _08880_ (.A1(_03257_),
    .A2(_03258_),
    .B1(_03259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03260_));
 sky130_fd_sc_hd__nor3_2 _08881_ (.A(_03257_),
    .B(_03258_),
    .C(_03259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03261_));
 sky130_fd_sc_hd__nor2_1 _08882_ (.A(_03260_),
    .B(_03261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03262_));
 sky130_fd_sc_hd__xnor2_1 _08883_ (.A(_03256_),
    .B(_03262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03263_));
 sky130_fd_sc_hd__xnor2_1 _08884_ (.A(_03250_),
    .B(_03263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03264_));
 sky130_fd_sc_hd__o21ba_1 _08885_ (.A1(_03234_),
    .A2(_03237_),
    .B1_N(_03235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03265_));
 sky130_fd_sc_hd__xnor2_1 _08886_ (.A(_03264_),
    .B(_03265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03266_));
 sky130_fd_sc_hd__a21oi_1 _08887_ (.A1(_03242_),
    .A2(_03243_),
    .B1(_03241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03267_));
 sky130_fd_sc_hd__xnor2_1 _08888_ (.A(_03266_),
    .B(_03267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03268_));
 sky130_fd_sc_hd__xnor2_1 _08889_ (.A(_03245_),
    .B(_03268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03269_));
 sky130_fd_sc_hd__xnor2_1 _08890_ (.A(_03207_),
    .B(_03269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03270_));
 sky130_fd_sc_hd__clkbuf_2 _08891_ (.A(_03193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03271_));
 sky130_fd_sc_hd__mux2_1 _08892_ (.A0(_03248_),
    .A1(_03270_),
    .S(_03271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03272_));
 sky130_fd_sc_hd__clkbuf_1 _08893_ (.A(_03272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[5] ));
 sky130_fd_sc_hd__nand2_1 _08894_ (.A(_03232_),
    .B(_03255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03273_));
 sky130_fd_sc_hd__or3_1 _08895_ (.A(_03256_),
    .B(_03260_),
    .C(_03261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03274_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08896_ (.A(\sa_inst.sak._03_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03275_));
 sky130_fd_sc_hd__a22oi_1 _08897_ (.A1(\sa_inst.sak._13_[6] ),
    .A2(_03229_),
    .B1(_03275_),
    .B2(\sa_inst.sak._13_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03276_));
 sky130_fd_sc_hd__and4_1 _08898_ (.A(\sa_inst.sak._13_[5] ),
    .B(\sa_inst.sak._13_[6] ),
    .C(_03229_),
    .D(\sa_inst.sak._03_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03277_));
 sky130_fd_sc_hd__nor2_1 _08899_ (.A(_03276_),
    .B(_03277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03278_));
 sky130_fd_sc_hd__nand2_1 _08900_ (.A(\sa_inst.sak._03_[7] ),
    .B(\sa_inst.sak._13_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03279_));
 sky130_fd_sc_hd__xnor2_1 _08901_ (.A(_03278_),
    .B(_03279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03280_));
 sky130_fd_sc_hd__or2_1 _08902_ (.A(_03252_),
    .B(_03254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03281_));
 sky130_fd_sc_hd__xor2_1 _08903_ (.A(_03280_),
    .B(_03281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03282_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08904_ (.A(\sa_inst.sak._13_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03283_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08905_ (.A(\sa_inst.sak._13_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03284_));
 sky130_fd_sc_hd__a22oi_1 _08906_ (.A1(_03196_),
    .A2(_03283_),
    .B1(_03284_),
    .B2(_03186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03285_));
 sky130_fd_sc_hd__and4_1 _08907_ (.A(_03186_),
    .B(_03213_),
    .C(\sa_inst.sak._13_[8] ),
    .D(\sa_inst.sak._13_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03286_));
 sky130_fd_sc_hd__nor2_1 _08908_ (.A(_03285_),
    .B(_03286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03287_));
 sky130_fd_sc_hd__xnor2_1 _08909_ (.A(_03282_),
    .B(_03287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03288_));
 sky130_fd_sc_hd__a21o_2 _08910_ (.A1(_03273_),
    .A2(_03274_),
    .B1(_03288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03289_));
 sky130_fd_sc_hd__nand3_1 _08911_ (.A(_03273_),
    .B(_03274_),
    .C(_03288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03290_));
 sky130_fd_sc_hd__o211ai_4 _08912_ (.A1(_03258_),
    .A2(_03261_),
    .B1(_03289_),
    .C1(_03290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03291_));
 sky130_fd_sc_hd__a211o_1 _08913_ (.A1(_03289_),
    .A2(_03290_),
    .B1(_03258_),
    .C1(_03261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03292_));
 sky130_fd_sc_hd__nand2_1 _08914_ (.A(_03250_),
    .B(_03263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03293_));
 sky130_fd_sc_hd__o21ai_1 _08915_ (.A1(_03264_),
    .A2(_03265_),
    .B1(_03293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03294_));
 sky130_fd_sc_hd__and3_1 _08916_ (.A(_03291_),
    .B(_03292_),
    .C(_03294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03295_));
 sky130_fd_sc_hd__a21oi_1 _08917_ (.A1(_03291_),
    .A2(_03292_),
    .B1(_03294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03296_));
 sky130_fd_sc_hd__or2_1 _08918_ (.A(_03295_),
    .B(_03296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03297_));
 sky130_fd_sc_hd__nor2_1 _08919_ (.A(_03266_),
    .B(_03267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03298_));
 sky130_fd_sc_hd__o21bai_1 _08920_ (.A1(_03245_),
    .A2(_03268_),
    .B1_N(_03298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03299_));
 sky130_fd_sc_hd__and2b_1 _08921_ (.A_N(_03297_),
    .B(_03299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03300_));
 sky130_fd_sc_hd__and2b_1 _08922_ (.A_N(_03299_),
    .B(_03297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03301_));
 sky130_fd_sc_hd__or2_1 _08923_ (.A(_03300_),
    .B(_03301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03302_));
 sky130_fd_sc_hd__xnor2_1 _08924_ (.A(_03207_),
    .B(_03302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03303_));
 sky130_fd_sc_hd__mux2_1 _08925_ (.A0(_03270_),
    .A1(_03303_),
    .S(_03271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03304_));
 sky130_fd_sc_hd__clkbuf_1 _08926_ (.A(_03304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[6] ));
 sky130_fd_sc_hd__nand2_1 _08927_ (.A(_03196_),
    .B(_03284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03305_));
 sky130_fd_sc_hd__a22oi_1 _08928_ (.A1(_03212_),
    .A2(_03230_),
    .B1(_03275_),
    .B2(_03201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03306_));
 sky130_fd_sc_hd__and4_1 _08929_ (.A(_03201_),
    .B(_03211_),
    .C(_03229_),
    .D(_03275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03307_));
 sky130_fd_sc_hd__nor2_1 _08930_ (.A(_03306_),
    .B(_03307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03308_));
 sky130_fd_sc_hd__nand2_1 _08931_ (.A(_03209_),
    .B(_03283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03309_));
 sky130_fd_sc_hd__xnor2_1 _08932_ (.A(_03308_),
    .B(_03309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03310_));
 sky130_fd_sc_hd__o21ba_1 _08933_ (.A1(_03276_),
    .A2(_03279_),
    .B1_N(_03277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03311_));
 sky130_fd_sc_hd__xnor2_1 _08934_ (.A(_03310_),
    .B(_03311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03312_));
 sky130_fd_sc_hd__xor2_1 _08935_ (.A(_03305_),
    .B(_03312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03313_));
 sky130_fd_sc_hd__a22o_1 _08936_ (.A1(_03280_),
    .A2(_03281_),
    .B1(_03282_),
    .B2(_03287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03314_));
 sky130_fd_sc_hd__xnor2_1 _08937_ (.A(_03313_),
    .B(_03314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03315_));
 sky130_fd_sc_hd__xnor2_1 _08938_ (.A(_03286_),
    .B(_03315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03316_));
 sky130_fd_sc_hd__nand2_1 _08939_ (.A(_03289_),
    .B(_03291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03317_));
 sky130_fd_sc_hd__xnor2_1 _08940_ (.A(_03316_),
    .B(_03317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03318_));
 sky130_fd_sc_hd__or3_1 _08941_ (.A(_03295_),
    .B(_03300_),
    .C(_03318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03319_));
 sky130_fd_sc_hd__o21ai_2 _08942_ (.A1(_03295_),
    .A2(_03300_),
    .B1(_03318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03320_));
 sky130_fd_sc_hd__nand2_1 _08943_ (.A(_03319_),
    .B(_03320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03321_));
 sky130_fd_sc_hd__xnor2_1 _08944_ (.A(_03207_),
    .B(_03321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03322_));
 sky130_fd_sc_hd__mux2_1 _08945_ (.A0(_03303_),
    .A1(_03322_),
    .S(_03271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03323_));
 sky130_fd_sc_hd__clkbuf_1 _08946_ (.A(_03323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[7] ));
 sky130_fd_sc_hd__a21o_1 _08947_ (.A1(_03289_),
    .A2(_03291_),
    .B1(_03316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03324_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08948_ (.A(_03275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03325_));
 sky130_fd_sc_hd__and2_1 _08949_ (.A(_03230_),
    .B(_03283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03326_));
 sky130_fd_sc_hd__a21oi_1 _08950_ (.A1(_03212_),
    .A2(_03325_),
    .B1(_03326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03327_));
 sky130_fd_sc_hd__and3_1 _08951_ (.A(_03212_),
    .B(_03275_),
    .C(_03326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03328_));
 sky130_fd_sc_hd__nor2_1 _08952_ (.A(_03327_),
    .B(_03328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03329_));
 sky130_fd_sc_hd__nand2_1 _08953_ (.A(_03209_),
    .B(_03284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03330_));
 sky130_fd_sc_hd__xnor2_1 _08954_ (.A(_03329_),
    .B(_03330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03331_));
 sky130_fd_sc_hd__o21ba_1 _08955_ (.A1(_03306_),
    .A2(_03309_),
    .B1_N(_03307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03332_));
 sky130_fd_sc_hd__inv_2 _08956_ (.A(_03332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03333_));
 sky130_fd_sc_hd__xnor2_1 _08957_ (.A(_03331_),
    .B(_03333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03334_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08958_ (.A(_03284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03335_));
 sky130_fd_sc_hd__and2b_1 _08959_ (.A_N(_03311_),
    .B(_03310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03336_));
 sky130_fd_sc_hd__a31oi_1 _08960_ (.A1(_03196_),
    .A2(_03335_),
    .A3(_03312_),
    .B1(_03336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03337_));
 sky130_fd_sc_hd__nor2_1 _08961_ (.A(_03334_),
    .B(_03337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03338_));
 sky130_fd_sc_hd__and2_1 _08962_ (.A(_03334_),
    .B(_03337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03339_));
 sky130_fd_sc_hd__and2b_1 _08963_ (.A_N(_03313_),
    .B(_03314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03340_));
 sky130_fd_sc_hd__a21oi_1 _08964_ (.A1(_03286_),
    .A2(_03315_),
    .B1(_03340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03341_));
 sky130_fd_sc_hd__or3_1 _08965_ (.A(_03338_),
    .B(_03339_),
    .C(_03341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03342_));
 sky130_fd_sc_hd__nor2_1 _08966_ (.A(_03338_),
    .B(_03339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03343_));
 sky130_fd_sc_hd__or2b_1 _08967_ (.A(_03343_),
    .B_N(_03341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03344_));
 sky130_fd_sc_hd__nand2_1 _08968_ (.A(_03342_),
    .B(_03344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03345_));
 sky130_fd_sc_hd__a21oi_1 _08969_ (.A1(_03324_),
    .A2(_03320_),
    .B1(_03345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03346_));
 sky130_fd_sc_hd__and3_1 _08970_ (.A(_03324_),
    .B(_03320_),
    .C(_03345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03347_));
 sky130_fd_sc_hd__nor2_1 _08971_ (.A(_03346_),
    .B(_03347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03348_));
 sky130_fd_sc_hd__xor2_1 _08972_ (.A(_02841_),
    .B(_03348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03349_));
 sky130_fd_sc_hd__mux2_1 _08973_ (.A0(_03322_),
    .A1(_03349_),
    .S(_03271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03350_));
 sky130_fd_sc_hd__clkbuf_1 _08974_ (.A(_03350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[8] ));
 sky130_fd_sc_hd__a21o_1 _08975_ (.A1(_03324_),
    .A2(_03320_),
    .B1(_03345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03351_));
 sky130_fd_sc_hd__a31o_1 _08976_ (.A1(_03209_),
    .A2(_03335_),
    .A3(_03329_),
    .B1(_03328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03352_));
 sky130_fd_sc_hd__a22oi_1 _08977_ (.A1(_03283_),
    .A2(_03325_),
    .B1(_03335_),
    .B2(_03230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03353_));
 sky130_fd_sc_hd__and4_1 _08978_ (.A(_03230_),
    .B(_03283_),
    .C(_03325_),
    .D(_03284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03354_));
 sky130_fd_sc_hd__nor2_1 _08979_ (.A(_03353_),
    .B(_03354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03355_));
 sky130_fd_sc_hd__xnor2_1 _08980_ (.A(_03352_),
    .B(_03355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03356_));
 sky130_fd_sc_hd__a21oi_1 _08981_ (.A1(_03331_),
    .A2(_03333_),
    .B1(_03338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03357_));
 sky130_fd_sc_hd__xnor2_1 _08982_ (.A(_03356_),
    .B(_03357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03358_));
 sky130_fd_sc_hd__a21oi_1 _08983_ (.A1(_03342_),
    .A2(_03351_),
    .B1(_03358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03359_));
 sky130_fd_sc_hd__and3_1 _08984_ (.A(_03342_),
    .B(_03351_),
    .C(_03358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03360_));
 sky130_fd_sc_hd__or2_1 _08985_ (.A(_03359_),
    .B(_03360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03361_));
 sky130_fd_sc_hd__xnor2_1 _08986_ (.A(_02841_),
    .B(_03361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03362_));
 sky130_fd_sc_hd__mux2_1 _08987_ (.A0(_03349_),
    .A1(_03362_),
    .S(_03271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03363_));
 sky130_fd_sc_hd__clkbuf_1 _08988_ (.A(_03363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[9] ));
 sky130_fd_sc_hd__inv_2 _08989_ (.A(_03356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03364_));
 sky130_fd_sc_hd__a21o_1 _08990_ (.A1(_03338_),
    .A2(_03364_),
    .B1(_03359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03365_));
 sky130_fd_sc_hd__and3b_1 _08991_ (.A_N(_03326_),
    .B(_03335_),
    .C(_03325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03366_));
 sky130_fd_sc_hd__and2_1 _08992_ (.A(_03352_),
    .B(_03355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03367_));
 sky130_fd_sc_hd__and3_1 _08993_ (.A(_03331_),
    .B(_03333_),
    .C(_03364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03368_));
 sky130_fd_sc_hd__nor2_1 _08994_ (.A(_03367_),
    .B(_03368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03369_));
 sky130_fd_sc_hd__xnor2_1 _08995_ (.A(_03366_),
    .B(_03369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03370_));
 sky130_fd_sc_hd__xnor2_1 _08996_ (.A(_03365_),
    .B(_03370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03371_));
 sky130_fd_sc_hd__xnor2_1 _08997_ (.A(_02841_),
    .B(_03371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03372_));
 sky130_fd_sc_hd__mux2_1 _08998_ (.A0(_03362_),
    .A1(_03372_),
    .S(_03193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03373_));
 sky130_fd_sc_hd__clkbuf_1 _08999_ (.A(_03373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[10] ));
 sky130_fd_sc_hd__a22o_1 _09000_ (.A1(_03366_),
    .A2(_03368_),
    .B1(_03370_),
    .B2(_03365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03374_));
 sky130_fd_sc_hd__o211a_1 _09001_ (.A1(_03326_),
    .A2(_03367_),
    .B1(_03325_),
    .C1(_03335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03375_));
 sky130_fd_sc_hd__xnor2_1 _09002_ (.A(_02840_),
    .B(_03375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03376_));
 sky130_fd_sc_hd__xnor2_1 _09003_ (.A(_03374_),
    .B(_03376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03377_));
 sky130_fd_sc_hd__mux2_1 _09004_ (.A0(_03372_),
    .A1(_03377_),
    .S(_03193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03378_));
 sky130_fd_sc_hd__clkbuf_1 _09005_ (.A(_03378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[11] ));
 sky130_fd_sc_hd__mux2_1 _09006_ (.A0(_03377_),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._01_ ),
    .S(_03193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03379_));
 sky130_fd_sc_hd__clkbuf_1 _09007_ (.A(_03379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[12] ));
 sky130_fd_sc_hd__buf_2 _09008_ (.A(\sa_inst.EOB_Q_o ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03380_));
 sky130_fd_sc_hd__clkbuf_2 _09009_ (.A(_03380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03381_));
 sky130_fd_sc_hd__mux2_1 _09010_ (.A0(\sa_inst.sak._06_[0] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[0] ),
    .S(_03381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03382_));
 sky130_fd_sc_hd__clkbuf_1 _09011_ (.A(_03382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ));
 sky130_fd_sc_hd__mux2_1 _09012_ (.A0(\sa_inst.sak._06_[1] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[1] ),
    .S(_03381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03383_));
 sky130_fd_sc_hd__clkbuf_1 _09013_ (.A(_03383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ));
 sky130_fd_sc_hd__mux2_1 _09014_ (.A0(\sa_inst.sak._06_[2] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[2] ),
    .S(_03381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03384_));
 sky130_fd_sc_hd__clkbuf_1 _09015_ (.A(_03384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ));
 sky130_fd_sc_hd__mux2_1 _09016_ (.A0(\sa_inst.sak._06_[3] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[3] ),
    .S(_03381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03385_));
 sky130_fd_sc_hd__clkbuf_1 _09017_ (.A(_03385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ));
 sky130_fd_sc_hd__mux2_1 _09018_ (.A0(\sa_inst.sak._06_[4] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[4] ),
    .S(_03381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03386_));
 sky130_fd_sc_hd__clkbuf_1 _09019_ (.A(_03386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ));
 sky130_fd_sc_hd__clkbuf_2 _09020_ (.A(_03380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03387_));
 sky130_fd_sc_hd__mux2_1 _09021_ (.A0(\sa_inst.sak._06_[5] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[5] ),
    .S(_03387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03388_));
 sky130_fd_sc_hd__clkbuf_1 _09022_ (.A(_03388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ));
 sky130_fd_sc_hd__mux2_1 _09023_ (.A0(\sa_inst.sak._06_[6] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[6] ),
    .S(_03387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03389_));
 sky130_fd_sc_hd__clkbuf_1 _09024_ (.A(_03389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ));
 sky130_fd_sc_hd__mux2_1 _09025_ (.A0(\sa_inst.sak._06_[7] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[7] ),
    .S(_03387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03390_));
 sky130_fd_sc_hd__clkbuf_1 _09026_ (.A(_03390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ));
 sky130_fd_sc_hd__mux2_1 _09027_ (.A0(\sa_inst.sak._06_[8] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[8] ),
    .S(_03387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03391_));
 sky130_fd_sc_hd__clkbuf_1 _09028_ (.A(_03391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ));
 sky130_fd_sc_hd__mux2_1 _09029_ (.A0(\sa_inst.sak._06_[9] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[9] ),
    .S(_03387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03392_));
 sky130_fd_sc_hd__clkbuf_1 _09030_ (.A(_03392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ));
 sky130_fd_sc_hd__clkbuf_2 _09031_ (.A(_03380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03393_));
 sky130_fd_sc_hd__mux2_1 _09032_ (.A0(\sa_inst.sak._06_[10] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[10] ),
    .S(_03393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03394_));
 sky130_fd_sc_hd__clkbuf_1 _09033_ (.A(_03394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ));
 sky130_fd_sc_hd__mux2_1 _09034_ (.A0(\sa_inst.sak._06_[11] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[11] ),
    .S(_03393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03395_));
 sky130_fd_sc_hd__clkbuf_1 _09035_ (.A(_03395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ));
 sky130_fd_sc_hd__mux2_1 _09036_ (.A0(\sa_inst.sak._06_[12] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[12] ),
    .S(_03393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03396_));
 sky130_fd_sc_hd__clkbuf_1 _09037_ (.A(_03396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ));
 sky130_fd_sc_hd__mux2_1 _09038_ (.A0(\sa_inst.sak._06_[13] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[13] ),
    .S(_03393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03397_));
 sky130_fd_sc_hd__clkbuf_1 _09039_ (.A(_03397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ));
 sky130_fd_sc_hd__mux2_1 _09040_ (.A0(\sa_inst.sak._06_[14] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[14] ),
    .S(_03393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03398_));
 sky130_fd_sc_hd__clkbuf_1 _09041_ (.A(_03398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ));
 sky130_fd_sc_hd__clkbuf_2 _09042_ (.A(_03380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03399_));
 sky130_fd_sc_hd__mux2_1 _09043_ (.A0(\sa_inst.sak._06_[15] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[15] ),
    .S(_03399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03400_));
 sky130_fd_sc_hd__clkbuf_1 _09044_ (.A(_03400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ));
 sky130_fd_sc_hd__mux2_1 _09045_ (.A0(\sa_inst.sak._06_[16] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[16] ),
    .S(_03399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03401_));
 sky130_fd_sc_hd__clkbuf_1 _09046_ (.A(_03401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ));
 sky130_fd_sc_hd__mux2_1 _09047_ (.A0(\sa_inst.sak._06_[17] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[17] ),
    .S(_03399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03402_));
 sky130_fd_sc_hd__clkbuf_1 _09048_ (.A(_03402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ));
 sky130_fd_sc_hd__mux2_1 _09049_ (.A0(\sa_inst.sak._06_[18] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[18] ),
    .S(_03399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03403_));
 sky130_fd_sc_hd__clkbuf_1 _09050_ (.A(_03403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ));
 sky130_fd_sc_hd__mux2_1 _09051_ (.A0(\sa_inst.sak._06_[19] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[19] ),
    .S(_03399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03404_));
 sky130_fd_sc_hd__clkbuf_1 _09052_ (.A(_03404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ));
 sky130_fd_sc_hd__buf_2 _09053_ (.A(\sa_inst.EOB_Q_o ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03405_));
 sky130_fd_sc_hd__buf_2 _09054_ (.A(_03405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03406_));
 sky130_fd_sc_hd__clkbuf_2 _09055_ (.A(_03406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03407_));
 sky130_fd_sc_hd__mux2_1 _09056_ (.A0(\sa_inst.sak._06_[20] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[20] ),
    .S(_03407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03408_));
 sky130_fd_sc_hd__clkbuf_1 _09057_ (.A(_03408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ));
 sky130_fd_sc_hd__mux2_1 _09058_ (.A0(\sa_inst.sak._06_[21] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[21] ),
    .S(_03407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03409_));
 sky130_fd_sc_hd__clkbuf_1 _09059_ (.A(_03409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ));
 sky130_fd_sc_hd__mux2_1 _09060_ (.A0(\sa_inst.sak._06_[22] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[22] ),
    .S(_03407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03410_));
 sky130_fd_sc_hd__clkbuf_1 _09061_ (.A(_03410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ));
 sky130_fd_sc_hd__mux2_1 _09062_ (.A0(\sa_inst.sak._06_[23] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[23] ),
    .S(_03407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03411_));
 sky130_fd_sc_hd__clkbuf_1 _09063_ (.A(_03411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ));
 sky130_fd_sc_hd__mux2_1 _09064_ (.A0(\sa_inst.sak._06_[24] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[24] ),
    .S(_03407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03412_));
 sky130_fd_sc_hd__clkbuf_1 _09065_ (.A(_03412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ));
 sky130_fd_sc_hd__clkbuf_2 _09066_ (.A(_03406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03413_));
 sky130_fd_sc_hd__mux2_1 _09067_ (.A0(\sa_inst.sak._06_[25] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[25] ),
    .S(_03413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03414_));
 sky130_fd_sc_hd__clkbuf_1 _09068_ (.A(_03414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ));
 sky130_fd_sc_hd__mux2_1 _09069_ (.A0(\sa_inst.sak._06_[26] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[26] ),
    .S(_03413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03415_));
 sky130_fd_sc_hd__clkbuf_1 _09070_ (.A(_03415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ));
 sky130_fd_sc_hd__mux2_1 _09071_ (.A0(\sa_inst.sak._06_[27] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[27] ),
    .S(_03413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03416_));
 sky130_fd_sc_hd__clkbuf_1 _09072_ (.A(_03416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ));
 sky130_fd_sc_hd__mux2_1 _09073_ (.A0(\sa_inst.sak._06_[28] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[28] ),
    .S(_03413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03417_));
 sky130_fd_sc_hd__clkbuf_1 _09074_ (.A(_03417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ));
 sky130_fd_sc_hd__mux2_1 _09075_ (.A0(\sa_inst.sak._06_[29] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[29] ),
    .S(_03413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03418_));
 sky130_fd_sc_hd__clkbuf_1 _09076_ (.A(_03418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ));
 sky130_fd_sc_hd__clkbuf_4 _09077_ (.A(_03406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03419_));
 sky130_fd_sc_hd__mux2_1 _09078_ (.A0(\sa_inst.sak._06_[30] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[30] ),
    .S(_03419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03420_));
 sky130_fd_sc_hd__clkbuf_1 _09079_ (.A(_03420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ));
 sky130_fd_sc_hd__mux2_1 _09080_ (.A0(\sa_inst.sak._06_[31] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[31] ),
    .S(_03419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03421_));
 sky130_fd_sc_hd__clkbuf_1 _09081_ (.A(_03421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ));
 sky130_fd_sc_hd__mux2_1 _09082_ (.A0(\sa_inst.sak._06_[32] ),
    .A1(\sa_inst.sak.rows:2.cols:3.pe_ij._02_ ),
    .S(_03419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03422_));
 sky130_fd_sc_hd__clkbuf_1 _09083_ (.A(_03422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ));
 sky130_fd_sc_hd__nand2_1 _09084_ (.A(_02766_),
    .B(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03423_));
 sky130_fd_sc_hd__xnor2_1 _09085_ (.A(_01824_),
    .B(_03423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[0] ));
 sky130_fd_sc_hd__and3_1 _09086_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[1] ),
    .B(_01839_),
    .C(_01842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03424_));
 sky130_fd_sc_hd__a21oi_1 _09087_ (.A1(_01840_),
    .A2(_01842_),
    .B1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03425_));
 sky130_fd_sc_hd__nand2_1 _09088_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[0] ),
    .B(_01824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03426_));
 sky130_fd_sc_hd__or3_1 _09089_ (.A(_03424_),
    .B(_03425_),
    .C(_03426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03427_));
 sky130_fd_sc_hd__o21ai_1 _09090_ (.A1(_03424_),
    .A2(_03425_),
    .B1(_03426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03428_));
 sky130_fd_sc_hd__a31o_1 _09091_ (.A1(_02132_),
    .A2(_03427_),
    .A3(_03428_),
    .B1(_01851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[1] ));
 sky130_fd_sc_hd__o21ba_1 _09092_ (.A1(_03425_),
    .A2(_03426_),
    .B1_N(_03424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03429_));
 sky130_fd_sc_hd__nor2_1 _09093_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[2] ),
    .B(_01861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03430_));
 sky130_fd_sc_hd__and2_1 _09094_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[2] ),
    .B(_01863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03431_));
 sky130_fd_sc_hd__or3_1 _09095_ (.A(_03429_),
    .B(_03430_),
    .C(_03431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03432_));
 sky130_fd_sc_hd__o21ai_1 _09096_ (.A1(_03430_),
    .A2(_03431_),
    .B1(_03429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03433_));
 sky130_fd_sc_hd__a31o_1 _09097_ (.A1(_02132_),
    .A2(_03432_),
    .A3(_03433_),
    .B1(_01868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[2] ));
 sky130_fd_sc_hd__nor2_1 _09098_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[3] ),
    .B(_01876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03434_));
 sky130_fd_sc_hd__or3b_1 _09099_ (.A(_01873_),
    .B(_01875_),
    .C_N(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03435_));
 sky130_fd_sc_hd__or2b_1 _09100_ (.A(_03434_),
    .B_N(_03435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03436_));
 sky130_fd_sc_hd__nand2_1 _09101_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[2] ),
    .B(_01863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03437_));
 sky130_fd_sc_hd__o21ai_1 _09102_ (.A1(_03429_),
    .A2(_03430_),
    .B1(_03437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03438_));
 sky130_fd_sc_hd__xnor2_1 _09103_ (.A(_03436_),
    .B(_03438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03439_));
 sky130_fd_sc_hd__mux2_1 _09104_ (.A0(_01876_),
    .A1(_03439_),
    .S(_02690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03440_));
 sky130_fd_sc_hd__clkbuf_1 _09105_ (.A(_03440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[3] ));
 sky130_fd_sc_hd__clkbuf_2 _09106_ (.A(_01883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03441_));
 sky130_fd_sc_hd__xnor2_1 _09107_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[4] ),
    .B(_01889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03442_));
 sky130_fd_sc_hd__o211a_1 _09108_ (.A1(_03429_),
    .A2(_03430_),
    .B1(_03437_),
    .C1(_03435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03443_));
 sky130_fd_sc_hd__or3_1 _09109_ (.A(_03434_),
    .B(_03442_),
    .C(_03443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03444_));
 sky130_fd_sc_hd__o21ai_1 _09110_ (.A1(_03434_),
    .A2(_03443_),
    .B1(_03442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03445_));
 sky130_fd_sc_hd__a31o_1 _09111_ (.A1(_03441_),
    .A2(_03444_),
    .A3(_03445_),
    .B1(_01894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[4] ));
 sky130_fd_sc_hd__xnor2_1 _09112_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[5] ),
    .B(_01899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03446_));
 sky130_fd_sc_hd__nand2_1 _09113_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[4] ),
    .B(_01889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03447_));
 sky130_fd_sc_hd__nand2_1 _09114_ (.A(_03447_),
    .B(_03444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03448_));
 sky130_fd_sc_hd__xnor2_1 _09115_ (.A(_03446_),
    .B(_03448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03449_));
 sky130_fd_sc_hd__mux2_1 _09116_ (.A0(_01900_),
    .A1(_03449_),
    .S(_02690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03450_));
 sky130_fd_sc_hd__clkbuf_1 _09117_ (.A(_03450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[5] ));
 sky130_fd_sc_hd__xnor2_1 _09118_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[6] ),
    .B(_01920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03451_));
 sky130_fd_sc_hd__nand2_1 _09119_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[5] ),
    .B(_01900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03452_));
 sky130_fd_sc_hd__nor2_1 _09120_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[5] ),
    .B(_01900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03453_));
 sky130_fd_sc_hd__a31o_1 _09121_ (.A1(_03447_),
    .A2(_03444_),
    .A3(_03452_),
    .B1(_03453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03454_));
 sky130_fd_sc_hd__or2_1 _09122_ (.A(_03451_),
    .B(_03454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03455_));
 sky130_fd_sc_hd__a21oi_1 _09123_ (.A1(_03451_),
    .A2(_03454_),
    .B1(_01924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03456_));
 sky130_fd_sc_hd__a22o_1 _09124_ (.A1(_02635_),
    .A2(_01921_),
    .B1(_03455_),
    .B2(_03456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[6] ));
 sky130_fd_sc_hd__buf_2 _09125_ (.A(_01978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03457_));
 sky130_fd_sc_hd__xnor2_1 _09126_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[7] ),
    .B(_01936_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03458_));
 sky130_fd_sc_hd__a21bo_1 _09127_ (.A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[6] ),
    .A2(_01921_),
    .B1_N(_03455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03459_));
 sky130_fd_sc_hd__xnor2_1 _09128_ (.A(_03458_),
    .B(_03459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03460_));
 sky130_fd_sc_hd__a21o_1 _09129_ (.A1(_03457_),
    .A2(_03460_),
    .B1(_01943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[7] ));
 sky130_fd_sc_hd__xnor2_1 _09130_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[8] ),
    .B(_01947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03461_));
 sky130_fd_sc_hd__o211a_1 _09131_ (.A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[7] ),
    .A2(_01936_),
    .B1(_01921_),
    .C1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03462_));
 sky130_fd_sc_hd__a21oi_1 _09132_ (.A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[7] ),
    .A2(_01936_),
    .B1(_03462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03463_));
 sky130_fd_sc_hd__a2111o_1 _09133_ (.A1(_03447_),
    .A2(_03452_),
    .B1(_03453_),
    .C1(_03451_),
    .D1(_03458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03464_));
 sky130_fd_sc_hd__or4_1 _09134_ (.A(_03444_),
    .B(_03446_),
    .C(_03451_),
    .D(_03458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03465_));
 sky130_fd_sc_hd__and3_1 _09135_ (.A(_03463_),
    .B(_03464_),
    .C(_03465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03466_));
 sky130_fd_sc_hd__a21o_1 _09136_ (.A1(_03461_),
    .A2(_03466_),
    .B1(_02093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03467_));
 sky130_fd_sc_hd__nor2_1 _09137_ (.A(_03461_),
    .B(_03466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03468_));
 sky130_fd_sc_hd__a2bb2o_1 _09138_ (.A1_N(_03467_),
    .A2_N(_03468_),
    .B1(_01948_),
    .B2(_01911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[8] ));
 sky130_fd_sc_hd__and3_1 _09139_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[9] ),
    .B(_01958_),
    .C(_01959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03469_));
 sky130_fd_sc_hd__nor2_1 _09140_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[9] ),
    .B(_01960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03470_));
 sky130_fd_sc_hd__a21oi_1 _09141_ (.A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[8] ),
    .A2(_01948_),
    .B1(_03468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03471_));
 sky130_fd_sc_hd__o21ai_1 _09142_ (.A1(_03469_),
    .A2(_03470_),
    .B1(_03471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03472_));
 sky130_fd_sc_hd__o31a_1 _09143_ (.A1(_03469_),
    .A2(_03470_),
    .A3(_03471_),
    .B1(_02766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03473_));
 sky130_fd_sc_hd__a22o_1 _09144_ (.A1(_02635_),
    .A2(_01960_),
    .B1(_03472_),
    .B2(_03473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[9] ));
 sky130_fd_sc_hd__xnor2_1 _09145_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[10] ),
    .B(_01976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03474_));
 sky130_fd_sc_hd__a21o_1 _09146_ (.A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[8] ),
    .A2(_01948_),
    .B1(_03469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03475_));
 sky130_fd_sc_hd__o21bai_1 _09147_ (.A1(_03468_),
    .A2(_03475_),
    .B1_N(_03470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03476_));
 sky130_fd_sc_hd__or2_1 _09148_ (.A(_03474_),
    .B(_03476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03477_));
 sky130_fd_sc_hd__nand2_1 _09149_ (.A(_03474_),
    .B(_03476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03478_));
 sky130_fd_sc_hd__a31o_1 _09150_ (.A1(_03441_),
    .A2(_03477_),
    .A3(_03478_),
    .B1(_01977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[10] ));
 sky130_fd_sc_hd__nand2_1 _09151_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[10] ),
    .B(_01976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03479_));
 sky130_fd_sc_hd__a21oi_1 _09152_ (.A1(_01982_),
    .A2(_01983_),
    .B1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03480_));
 sky130_fd_sc_hd__and3_1 _09153_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[11] ),
    .B(_01982_),
    .C(_01983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03481_));
 sky130_fd_sc_hd__or2_1 _09154_ (.A(_03480_),
    .B(_03481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03482_));
 sky130_fd_sc_hd__a21o_1 _09155_ (.A1(_03479_),
    .A2(_03477_),
    .B1(_03482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03483_));
 sky130_fd_sc_hd__nand3_1 _09156_ (.A(_03479_),
    .B(_03477_),
    .C(_03482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03484_));
 sky130_fd_sc_hd__a31o_1 _09157_ (.A1(_03441_),
    .A2(_03483_),
    .A3(_03484_),
    .B1(_01989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[11] ));
 sky130_fd_sc_hd__o21ba_1 _09158_ (.A1(_03479_),
    .A2(_03480_),
    .B1_N(_03481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03485_));
 sky130_fd_sc_hd__or3_1 _09159_ (.A(_03474_),
    .B(_03480_),
    .C(_03481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03486_));
 sky130_fd_sc_hd__or3b_1 _09160_ (.A(_03470_),
    .B(_03486_),
    .C_N(_03475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03487_));
 sky130_fd_sc_hd__or3_1 _09161_ (.A(_03461_),
    .B(_03469_),
    .C(_03470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03488_));
 sky130_fd_sc_hd__a311o_1 _09162_ (.A1(_03463_),
    .A2(_03464_),
    .A3(_03465_),
    .B1(_03488_),
    .C1(_03486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03489_));
 sky130_fd_sc_hd__nand2_1 _09163_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[12] ),
    .B(_02001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03490_));
 sky130_fd_sc_hd__or2_1 _09164_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[12] ),
    .B(_02000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03491_));
 sky130_fd_sc_hd__nand2_1 _09165_ (.A(_03490_),
    .B(_03491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03492_));
 sky130_fd_sc_hd__a31o_1 _09166_ (.A1(_03485_),
    .A2(_03487_),
    .A3(_03489_),
    .B1(_03492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03493_));
 sky130_fd_sc_hd__o211ai_1 _09167_ (.A1(_03476_),
    .A2(_03486_),
    .B1(_03485_),
    .C1(_03492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03494_));
 sky130_fd_sc_hd__a31o_1 _09168_ (.A1(_03441_),
    .A2(_03493_),
    .A3(_03494_),
    .B1(_02005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[12] ));
 sky130_fd_sc_hd__inv_2 _09169_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03495_));
 sky130_fd_sc_hd__nor2_1 _09170_ (.A(_03495_),
    .B(_02013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03496_));
 sky130_fd_sc_hd__and2_1 _09171_ (.A(_03495_),
    .B(_02013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03497_));
 sky130_fd_sc_hd__nor2_1 _09172_ (.A(_03496_),
    .B(_03497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03498_));
 sky130_fd_sc_hd__nand2_1 _09173_ (.A(_03490_),
    .B(_03493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03499_));
 sky130_fd_sc_hd__xor2_1 _09174_ (.A(_03498_),
    .B(_03499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03500_));
 sky130_fd_sc_hd__a21o_1 _09175_ (.A1(_03457_),
    .A2(_03500_),
    .B1(_02014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[13] ));
 sky130_fd_sc_hd__xnor2_1 _09176_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[14] ),
    .B(_02021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03501_));
 sky130_fd_sc_hd__or2_1 _09177_ (.A(_03495_),
    .B(_02013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03502_));
 sky130_fd_sc_hd__a31o_1 _09178_ (.A1(_03490_),
    .A2(_03493_),
    .A3(_03502_),
    .B1(_03497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03503_));
 sky130_fd_sc_hd__or2_1 _09179_ (.A(_03501_),
    .B(_03503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03504_));
 sky130_fd_sc_hd__nand2_1 _09180_ (.A(_03501_),
    .B(_03503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03505_));
 sky130_fd_sc_hd__a31o_1 _09181_ (.A1(_03441_),
    .A2(_03504_),
    .A3(_03505_),
    .B1(_02022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[14] ));
 sky130_fd_sc_hd__clkbuf_2 _09182_ (.A(_01883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03506_));
 sky130_fd_sc_hd__nand2_1 _09183_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[14] ),
    .B(_02021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03507_));
 sky130_fd_sc_hd__xnor2_1 _09184_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[15] ),
    .B(_02026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03508_));
 sky130_fd_sc_hd__a21o_1 _09185_ (.A1(_03507_),
    .A2(_03504_),
    .B1(_03508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03509_));
 sky130_fd_sc_hd__nand3_1 _09186_ (.A(_03507_),
    .B(_03504_),
    .C(_03508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03510_));
 sky130_fd_sc_hd__a31o_1 _09187_ (.A1(_03506_),
    .A2(_03509_),
    .A3(_03510_),
    .B1(_02031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[15] ));
 sky130_fd_sc_hd__nor2_1 _09188_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[15] ),
    .B(_02026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03511_));
 sky130_fd_sc_hd__nor2_1 _09189_ (.A(_03501_),
    .B(_03508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03512_));
 sky130_fd_sc_hd__nand2_1 _09190_ (.A(_03498_),
    .B(_03512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03513_));
 sky130_fd_sc_hd__o21ai_1 _09191_ (.A1(_03490_),
    .A2(_03497_),
    .B1(_03502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03514_));
 sky130_fd_sc_hd__a22oi_1 _09192_ (.A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[15] ),
    .A2(_02026_),
    .B1(_03512_),
    .B2(_03514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03515_));
 sky130_fd_sc_hd__o221a_2 _09193_ (.A1(_03507_),
    .A2(_03511_),
    .B1(_03513_),
    .B2(_03493_),
    .C1(_03515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03516_));
 sky130_fd_sc_hd__xnor2_1 _09194_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[16] ),
    .B(_02055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03517_));
 sky130_fd_sc_hd__nor2_1 _09195_ (.A(_03516_),
    .B(_03517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03518_));
 sky130_fd_sc_hd__a21o_1 _09196_ (.A1(_03516_),
    .A2(_03517_),
    .B1(_02093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03519_));
 sky130_fd_sc_hd__o21bai_1 _09197_ (.A1(_03518_),
    .A2(_03519_),
    .B1_N(_02095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[16] ));
 sky130_fd_sc_hd__a21oi_1 _09198_ (.A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[16] ),
    .A2(_02046_),
    .B1(_03518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03520_));
 sky130_fd_sc_hd__nand2_1 _09199_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[17] ),
    .B(_02055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03521_));
 sky130_fd_sc_hd__or2_1 _09200_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[17] ),
    .B(_02037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03522_));
 sky130_fd_sc_hd__nand2_1 _09201_ (.A(_03521_),
    .B(_03522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03523_));
 sky130_fd_sc_hd__or2_1 _09202_ (.A(_03520_),
    .B(_03523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03524_));
 sky130_fd_sc_hd__nand2_1 _09203_ (.A(_03520_),
    .B(_03523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03525_));
 sky130_fd_sc_hd__a31o_1 _09204_ (.A1(_03506_),
    .A2(_03524_),
    .A3(_03525_),
    .B1(_02137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[17] ));
 sky130_fd_sc_hd__or2b_1 _09205_ (.A(_03520_),
    .B_N(_03522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03526_));
 sky130_fd_sc_hd__nand2_1 _09206_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[18] ),
    .B(_02055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03527_));
 sky130_fd_sc_hd__or2_1 _09207_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[18] ),
    .B(_02037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03528_));
 sky130_fd_sc_hd__nand2_1 _09208_ (.A(_03527_),
    .B(_03528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03529_));
 sky130_fd_sc_hd__a21o_1 _09209_ (.A1(_03521_),
    .A2(_03526_),
    .B1(_03529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03530_));
 sky130_fd_sc_hd__nand3_1 _09210_ (.A(_03521_),
    .B(_03526_),
    .C(_03529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03531_));
 sky130_fd_sc_hd__a31o_1 _09211_ (.A1(_03506_),
    .A2(_03530_),
    .A3(_03531_),
    .B1(_02137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[18] ));
 sky130_fd_sc_hd__xnor2_1 _09212_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[19] ),
    .B(_02041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03532_));
 sky130_fd_sc_hd__a21o_1 _09213_ (.A1(_03527_),
    .A2(_03530_),
    .B1(_03532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03533_));
 sky130_fd_sc_hd__nand3_1 _09214_ (.A(_03527_),
    .B(_03530_),
    .C(_03532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03534_));
 sky130_fd_sc_hd__clkbuf_2 _09215_ (.A(_02048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03535_));
 sky130_fd_sc_hd__a31o_1 _09216_ (.A1(_03506_),
    .A2(_03533_),
    .A3(_03534_),
    .B1(_03535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[19] ));
 sky130_fd_sc_hd__and2_1 _09217_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[20] ),
    .B(_02053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03536_));
 sky130_fd_sc_hd__nor2_1 _09218_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[20] ),
    .B(_02042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03537_));
 sky130_fd_sc_hd__or2_1 _09219_ (.A(_03536_),
    .B(_03537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03538_));
 sky130_fd_sc_hd__or4_1 _09220_ (.A(_03517_),
    .B(_03523_),
    .C(_03529_),
    .D(_03532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03539_));
 sky130_fd_sc_hd__o41a_1 _09221_ (.A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[16] ),
    .A2(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[17] ),
    .A3(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[18] ),
    .A4(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[19] ),
    .B1(_02123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03540_));
 sky130_fd_sc_hd__o21ba_1 _09222_ (.A1(_03516_),
    .A2(_03539_),
    .B1_N(_03540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03541_));
 sky130_fd_sc_hd__nor2_1 _09223_ (.A(_03538_),
    .B(_03541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03542_));
 sky130_fd_sc_hd__a21o_1 _09224_ (.A1(_03538_),
    .A2(_03541_),
    .B1(_02093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03543_));
 sky130_fd_sc_hd__o21bai_1 _09225_ (.A1(_03542_),
    .A2(_03543_),
    .B1_N(_02095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[20] ));
 sky130_fd_sc_hd__or2_1 _09226_ (.A(_03536_),
    .B(_03542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03544_));
 sky130_fd_sc_hd__and2_1 _09227_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[21] ),
    .B(_02053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03545_));
 sky130_fd_sc_hd__or2_1 _09228_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[21] ),
    .B(_02053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03546_));
 sky130_fd_sc_hd__or2b_1 _09229_ (.A(_03545_),
    .B_N(_03546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03547_));
 sky130_fd_sc_hd__xnor2_1 _09230_ (.A(_03544_),
    .B(_03547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03548_));
 sky130_fd_sc_hd__a21o_1 _09231_ (.A1(_03457_),
    .A2(_03548_),
    .B1(_02050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[21] ));
 sky130_fd_sc_hd__xor2_1 _09232_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[22] ),
    .B(_02042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03549_));
 sky130_fd_sc_hd__o311a_1 _09233_ (.A1(_03536_),
    .A2(_03542_),
    .A3(_03545_),
    .B1(_03546_),
    .C1(_03549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03550_));
 sky130_fd_sc_hd__inv_2 _09234_ (.A(_03550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03551_));
 sky130_fd_sc_hd__a211o_1 _09235_ (.A1(_03544_),
    .A2(_03546_),
    .B1(_03549_),
    .C1(_03545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03552_));
 sky130_fd_sc_hd__a31o_1 _09236_ (.A1(_03506_),
    .A2(_03551_),
    .A3(_03552_),
    .B1(_03535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[22] ));
 sky130_fd_sc_hd__xor2_1 _09237_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[23] ),
    .B(_02042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03553_));
 sky130_fd_sc_hd__a21oi_1 _09238_ (.A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[22] ),
    .A2(_02107_),
    .B1(_03550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03554_));
 sky130_fd_sc_hd__xnor2_1 _09239_ (.A(_03553_),
    .B(_03554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03555_));
 sky130_fd_sc_hd__a21o_1 _09240_ (.A1(_03457_),
    .A2(_03555_),
    .B1(_02060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[23] ));
 sky130_fd_sc_hd__nand2_1 _09241_ (.A(_03549_),
    .B(_03553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03556_));
 sky130_fd_sc_hd__or4_1 _09242_ (.A(_03538_),
    .B(_03539_),
    .C(_03547_),
    .D(_03556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03557_));
 sky130_fd_sc_hd__o41a_1 _09243_ (.A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[20] ),
    .A2(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[21] ),
    .A3(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[22] ),
    .A4(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[23] ),
    .B1(_02123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03558_));
 sky130_fd_sc_hd__nor2_1 _09244_ (.A(_03540_),
    .B(_03558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03559_));
 sky130_fd_sc_hd__o21ai_4 _09245_ (.A1(_03516_),
    .A2(_03557_),
    .B1(_03559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03560_));
 sky130_fd_sc_hd__xor2_1 _09246_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[24] ),
    .B(_02123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03561_));
 sky130_fd_sc_hd__nand2_1 _09247_ (.A(_03560_),
    .B(_03561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03562_));
 sky130_fd_sc_hd__or2_1 _09248_ (.A(_03560_),
    .B(_03561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03563_));
 sky130_fd_sc_hd__a31o_1 _09249_ (.A1(_02691_),
    .A2(_03562_),
    .A3(_03563_),
    .B1(_03535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[24] ));
 sky130_fd_sc_hd__xor2_1 _09250_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[25] ),
    .B(_02123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03564_));
 sky130_fd_sc_hd__a22o_1 _09251_ (.A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[24] ),
    .A2(_02107_),
    .B1(_03560_),
    .B2(_03561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03565_));
 sky130_fd_sc_hd__xor2_1 _09252_ (.A(_03564_),
    .B(_03565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03566_));
 sky130_fd_sc_hd__a21o_1 _09253_ (.A1(_03457_),
    .A2(_03566_),
    .B1(_02060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[25] ));
 sky130_fd_sc_hd__o21ai_1 _09254_ (.A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[24] ),
    .A2(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[25] ),
    .B1(_02110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03567_));
 sky130_fd_sc_hd__and2_1 _09255_ (.A(_03561_),
    .B(_03564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03568_));
 sky130_fd_sc_hd__nand2_1 _09256_ (.A(_03560_),
    .B(_03568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03569_));
 sky130_fd_sc_hd__nand2_1 _09257_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[26] ),
    .B(_02077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03570_));
 sky130_fd_sc_hd__or2_1 _09258_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[26] ),
    .B(_02043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03571_));
 sky130_fd_sc_hd__nand2_1 _09259_ (.A(_03570_),
    .B(_03571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03572_));
 sky130_fd_sc_hd__a21o_1 _09260_ (.A1(_03567_),
    .A2(_03569_),
    .B1(_03572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03573_));
 sky130_fd_sc_hd__nand3_1 _09261_ (.A(_03572_),
    .B(_03567_),
    .C(_03569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03574_));
 sky130_fd_sc_hd__a31o_1 _09262_ (.A1(_02691_),
    .A2(_03573_),
    .A3(_03574_),
    .B1(_03535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[26] ));
 sky130_fd_sc_hd__xnor2_1 _09263_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[27] ),
    .B(_02044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03575_));
 sky130_fd_sc_hd__nand2_1 _09264_ (.A(_03570_),
    .B(_03573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03576_));
 sky130_fd_sc_hd__xnor2_1 _09265_ (.A(_03575_),
    .B(_03576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03577_));
 sky130_fd_sc_hd__a21o_1 _09266_ (.A1(_01829_),
    .A2(_03577_),
    .B1(_02060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[27] ));
 sky130_fd_sc_hd__nor2_1 _09267_ (.A(_03572_),
    .B(_03575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03578_));
 sky130_fd_sc_hd__o41a_1 _09268_ (.A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[24] ),
    .A2(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[25] ),
    .A3(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[26] ),
    .A4(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[27] ),
    .B1(_02124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03579_));
 sky130_fd_sc_hd__a31oi_2 _09269_ (.A1(_03560_),
    .A2(_03568_),
    .A3(_03578_),
    .B1(_03579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03580_));
 sky130_fd_sc_hd__and2_1 _09270_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[28] ),
    .B(_02044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03581_));
 sky130_fd_sc_hd__nor2_1 _09271_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[28] ),
    .B(_02124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03582_));
 sky130_fd_sc_hd__or2_1 _09272_ (.A(_03581_),
    .B(_03582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03583_));
 sky130_fd_sc_hd__nor2_1 _09273_ (.A(_03580_),
    .B(_03583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03584_));
 sky130_fd_sc_hd__a21o_1 _09274_ (.A1(_03580_),
    .A2(_03583_),
    .B1(_02093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03585_));
 sky130_fd_sc_hd__o21bai_1 _09275_ (.A1(_03584_),
    .A2(_03585_),
    .B1_N(_02049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[28] ));
 sky130_fd_sc_hd__nand2_1 _09276_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[29] ),
    .B(_02045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03586_));
 sky130_fd_sc_hd__or2_1 _09277_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[29] ),
    .B(_02045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03587_));
 sky130_fd_sc_hd__o211ai_1 _09278_ (.A1(_03581_),
    .A2(_03584_),
    .B1(_03586_),
    .C1(_03587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03588_));
 sky130_fd_sc_hd__a211o_1 _09279_ (.A1(_03586_),
    .A2(_03587_),
    .B1(_03581_),
    .C1(_03584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03589_));
 sky130_fd_sc_hd__a31o_1 _09280_ (.A1(_02691_),
    .A2(_03588_),
    .A3(_03589_),
    .B1(_03535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[29] ));
 sky130_fd_sc_hd__o21ai_1 _09281_ (.A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[28] ),
    .A2(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[29] ),
    .B1(_02047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03590_));
 sky130_fd_sc_hd__or4bb_1 _09282_ (.A(_03580_),
    .B(_03583_),
    .C_N(_03586_),
    .D_N(_03587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03591_));
 sky130_fd_sc_hd__nand2_1 _09283_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[30] ),
    .B(_02110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03592_));
 sky130_fd_sc_hd__or2_1 _09284_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[30] ),
    .B(_02110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03593_));
 sky130_fd_sc_hd__nand2_1 _09285_ (.A(_03592_),
    .B(_03593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03594_));
 sky130_fd_sc_hd__a21o_1 _09286_ (.A1(_03590_),
    .A2(_03591_),
    .B1(_03594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03595_));
 sky130_fd_sc_hd__nand3_1 _09287_ (.A(_03594_),
    .B(_03590_),
    .C(_03591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03596_));
 sky130_fd_sc_hd__a31o_1 _09288_ (.A1(_02691_),
    .A2(_03595_),
    .A3(_03596_),
    .B1(_02095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[30] ));
 sky130_fd_sc_hd__xnor2_1 _09289_ (.A(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[31] ),
    .B(_02107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03597_));
 sky130_fd_sc_hd__a21oi_1 _09290_ (.A1(_03592_),
    .A2(_03595_),
    .B1(_03597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03598_));
 sky130_fd_sc_hd__a31o_1 _09291_ (.A1(_03592_),
    .A2(_03595_),
    .A3(_03597_),
    .B1(_01910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03599_));
 sky130_fd_sc_hd__o21bai_1 _09292_ (.A1(_03598_),
    .A2(_03599_),
    .B1_N(_02049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[31] ));
 sky130_fd_sc_hd__mux2_1 _09293_ (.A0(\sa_inst.sak._12_[0] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[0] ),
    .S(_02838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03600_));
 sky130_fd_sc_hd__clkbuf_1 _09294_ (.A(_03600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ));
 sky130_fd_sc_hd__mux2_1 _09295_ (.A0(\sa_inst.sak._12_[1] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[1] ),
    .S(_02838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03601_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09296_ (.A(_03601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ));
 sky130_fd_sc_hd__mux2_1 _09297_ (.A0(\sa_inst.sak._12_[2] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[2] ),
    .S(_02838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03602_));
 sky130_fd_sc_hd__clkbuf_1 _09298_ (.A(_03602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ));
 sky130_fd_sc_hd__mux2_1 _09299_ (.A0(\sa_inst.sak._12_[3] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[3] ),
    .S(_02838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03603_));
 sky130_fd_sc_hd__clkbuf_1 _09300_ (.A(_03603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ));
 sky130_fd_sc_hd__clkbuf_2 _09301_ (.A(_02831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03604_));
 sky130_fd_sc_hd__mux2_1 _09302_ (.A0(\sa_inst.sak._12_[4] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[4] ),
    .S(_03604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03605_));
 sky130_fd_sc_hd__clkbuf_1 _09303_ (.A(_03605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ));
 sky130_fd_sc_hd__mux2_1 _09304_ (.A0(\sa_inst.sak._12_[5] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[5] ),
    .S(_03604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03606_));
 sky130_fd_sc_hd__clkbuf_1 _09305_ (.A(_03606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ));
 sky130_fd_sc_hd__mux2_1 _09306_ (.A0(\sa_inst.sak._12_[6] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[6] ),
    .S(_03604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03607_));
 sky130_fd_sc_hd__clkbuf_1 _09307_ (.A(_03607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ));
 sky130_fd_sc_hd__mux2_1 _09308_ (.A0(\sa_inst.sak._12_[7] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[7] ),
    .S(_03604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03608_));
 sky130_fd_sc_hd__clkbuf_1 _09309_ (.A(_03608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ));
 sky130_fd_sc_hd__mux2_1 _09310_ (.A0(\sa_inst.sak._12_[8] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[8] ),
    .S(_03604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03609_));
 sky130_fd_sc_hd__clkbuf_1 _09311_ (.A(_03609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ));
 sky130_fd_sc_hd__clkbuf_2 _09312_ (.A(_02831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03610_));
 sky130_fd_sc_hd__mux2_1 _09313_ (.A0(\sa_inst.sak._12_[9] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[9] ),
    .S(_03610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03611_));
 sky130_fd_sc_hd__clkbuf_1 _09314_ (.A(_03611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ));
 sky130_fd_sc_hd__mux2_1 _09315_ (.A0(\sa_inst.sak._12_[10] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[10] ),
    .S(_03610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03612_));
 sky130_fd_sc_hd__clkbuf_1 _09316_ (.A(_03612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ));
 sky130_fd_sc_hd__mux2_1 _09317_ (.A0(\sa_inst.sak._12_[11] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[11] ),
    .S(_03610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03613_));
 sky130_fd_sc_hd__clkbuf_1 _09318_ (.A(_03613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ));
 sky130_fd_sc_hd__mux2_1 _09319_ (.A0(\sa_inst.sak._12_[12] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[12] ),
    .S(_03610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03614_));
 sky130_fd_sc_hd__clkbuf_1 _09320_ (.A(_03614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ));
 sky130_fd_sc_hd__mux2_1 _09321_ (.A0(\sa_inst.sak._12_[13] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[13] ),
    .S(_03610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03615_));
 sky130_fd_sc_hd__clkbuf_1 _09322_ (.A(_03615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ));
 sky130_fd_sc_hd__clkbuf_2 _09323_ (.A(_02831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03616_));
 sky130_fd_sc_hd__mux2_1 _09324_ (.A0(\sa_inst.sak._12_[14] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[14] ),
    .S(_03616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03617_));
 sky130_fd_sc_hd__clkbuf_1 _09325_ (.A(_03617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ));
 sky130_fd_sc_hd__mux2_1 _09326_ (.A0(\sa_inst.sak._12_[15] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[15] ),
    .S(_03616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03618_));
 sky130_fd_sc_hd__clkbuf_1 _09327_ (.A(_03618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ));
 sky130_fd_sc_hd__mux2_1 _09328_ (.A0(\sa_inst.sak._12_[16] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[16] ),
    .S(_03616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03619_));
 sky130_fd_sc_hd__clkbuf_1 _09329_ (.A(_03619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ));
 sky130_fd_sc_hd__mux2_1 _09330_ (.A0(\sa_inst.sak._12_[17] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[17] ),
    .S(_03616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03620_));
 sky130_fd_sc_hd__clkbuf_1 _09331_ (.A(_03620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ));
 sky130_fd_sc_hd__mux2_1 _09332_ (.A0(\sa_inst.sak._12_[18] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[18] ),
    .S(_03616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03621_));
 sky130_fd_sc_hd__clkbuf_1 _09333_ (.A(_03621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ));
 sky130_fd_sc_hd__clkbuf_2 _09334_ (.A(_02796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03622_));
 sky130_fd_sc_hd__mux2_1 _09335_ (.A0(\sa_inst.sak._12_[19] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[19] ),
    .S(_03622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03623_));
 sky130_fd_sc_hd__clkbuf_1 _09336_ (.A(_03623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ));
 sky130_fd_sc_hd__mux2_1 _09337_ (.A0(\sa_inst.sak._12_[20] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[20] ),
    .S(_03622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03624_));
 sky130_fd_sc_hd__clkbuf_1 _09338_ (.A(_03624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ));
 sky130_fd_sc_hd__mux2_1 _09339_ (.A0(\sa_inst.sak._12_[21] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[21] ),
    .S(_03622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03625_));
 sky130_fd_sc_hd__clkbuf_1 _09340_ (.A(_03625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ));
 sky130_fd_sc_hd__mux2_1 _09341_ (.A0(\sa_inst.sak._12_[22] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[22] ),
    .S(_03622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03626_));
 sky130_fd_sc_hd__clkbuf_1 _09342_ (.A(_03626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ));
 sky130_fd_sc_hd__mux2_1 _09343_ (.A0(\sa_inst.sak._12_[23] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[23] ),
    .S(_03622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03627_));
 sky130_fd_sc_hd__clkbuf_1 _09344_ (.A(_03627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ));
 sky130_fd_sc_hd__clkbuf_2 _09345_ (.A(_02796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03628_));
 sky130_fd_sc_hd__mux2_1 _09346_ (.A0(\sa_inst.sak._12_[24] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[24] ),
    .S(_03628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03629_));
 sky130_fd_sc_hd__clkbuf_1 _09347_ (.A(_03629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ));
 sky130_fd_sc_hd__mux2_1 _09348_ (.A0(\sa_inst.sak._12_[25] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[25] ),
    .S(_03628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03630_));
 sky130_fd_sc_hd__clkbuf_1 _09349_ (.A(_03630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ));
 sky130_fd_sc_hd__mux2_1 _09350_ (.A0(\sa_inst.sak._12_[26] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[26] ),
    .S(_03628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03631_));
 sky130_fd_sc_hd__clkbuf_1 _09351_ (.A(_03631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ));
 sky130_fd_sc_hd__mux2_1 _09352_ (.A0(\sa_inst.sak._12_[27] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[27] ),
    .S(_03628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03632_));
 sky130_fd_sc_hd__clkbuf_1 _09353_ (.A(_03632_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ));
 sky130_fd_sc_hd__mux2_1 _09354_ (.A0(\sa_inst.sak._12_[28] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[28] ),
    .S(_03628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03633_));
 sky130_fd_sc_hd__clkbuf_1 _09355_ (.A(_03633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ));
 sky130_fd_sc_hd__buf_4 _09356_ (.A(_02796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03634_));
 sky130_fd_sc_hd__mux2_1 _09357_ (.A0(\sa_inst.sak._12_[29] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[29] ),
    .S(_03634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03635_));
 sky130_fd_sc_hd__clkbuf_1 _09358_ (.A(_03635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ));
 sky130_fd_sc_hd__mux2_1 _09359_ (.A0(\sa_inst.sak._12_[30] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[30] ),
    .S(_03634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03636_));
 sky130_fd_sc_hd__clkbuf_1 _09360_ (.A(_03636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ));
 sky130_fd_sc_hd__mux2_1 _09361_ (.A0(\sa_inst.sak._12_[31] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[31] ),
    .S(_03634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03637_));
 sky130_fd_sc_hd__clkbuf_1 _09362_ (.A(_03637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ));
 sky130_fd_sc_hd__mux2_1 _09363_ (.A0(\sa_inst.sak._12_[32] ),
    .A1(\sa_inst.sak.rows:3.cols:1.pe_ij._02_ ),
    .S(_03634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03638_));
 sky130_fd_sc_hd__clkbuf_1 _09364_ (.A(_03638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ));
 sky130_fd_sc_hd__nand2_1 _09365_ (.A(_02854_),
    .B(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03639_));
 sky130_fd_sc_hd__xnor2_1 _09366_ (.A(_02852_),
    .B(_03639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[0] ));
 sky130_fd_sc_hd__and3_1 _09367_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[1] ),
    .B(_02866_),
    .C(_02868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03640_));
 sky130_fd_sc_hd__a21o_1 _09368_ (.A1(_02866_),
    .A2(_02868_),
    .B1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03641_));
 sky130_fd_sc_hd__or2b_1 _09369_ (.A(_03640_),
    .B_N(_03641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03642_));
 sky130_fd_sc_hd__nand2_1 _09370_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[0] ),
    .B(_02852_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03643_));
 sky130_fd_sc_hd__xor2_1 _09371_ (.A(_03642_),
    .B(_03643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03644_));
 sky130_fd_sc_hd__mux2_1 _09372_ (.A0(_02869_),
    .A1(_03644_),
    .S(_02914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03645_));
 sky130_fd_sc_hd__clkbuf_1 _09373_ (.A(_03645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[1] ));
 sky130_fd_sc_hd__a31o_1 _09374_ (.A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[0] ),
    .A2(_02852_),
    .A3(_03641_),
    .B1(_03640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03646_));
 sky130_fd_sc_hd__or2_1 _09375_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[2] ),
    .B(_02892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03647_));
 sky130_fd_sc_hd__nand2_1 _09376_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[2] ),
    .B(_02892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03648_));
 sky130_fd_sc_hd__nand3_1 _09377_ (.A(_03646_),
    .B(_03647_),
    .C(_03648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03649_));
 sky130_fd_sc_hd__a21o_1 _09378_ (.A1(_03647_),
    .A2(_03648_),
    .B1(_03646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03650_));
 sky130_fd_sc_hd__a31o_1 _09379_ (.A1(_03170_),
    .A2(_03649_),
    .A3(_03650_),
    .B1(_02899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[2] ));
 sky130_fd_sc_hd__or2_1 _09380_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[3] ),
    .B(_02907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03651_));
 sky130_fd_sc_hd__nand2_1 _09381_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[3] ),
    .B(_02907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03652_));
 sky130_fd_sc_hd__nand2_1 _09382_ (.A(_03651_),
    .B(_03652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03653_));
 sky130_fd_sc_hd__and2_1 _09383_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[2] ),
    .B(_02892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03654_));
 sky130_fd_sc_hd__a21o_1 _09384_ (.A1(_03646_),
    .A2(_03647_),
    .B1(_03654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03655_));
 sky130_fd_sc_hd__xnor2_1 _09385_ (.A(_03653_),
    .B(_03655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03656_));
 sky130_fd_sc_hd__mux2_1 _09386_ (.A0(_02907_),
    .A1(_03656_),
    .S(_02914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03657_));
 sky130_fd_sc_hd__clkbuf_1 _09387_ (.A(_03657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[3] ));
 sky130_fd_sc_hd__nor2_1 _09388_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[3] ),
    .B(_02907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03658_));
 sky130_fd_sc_hd__xnor2_1 _09389_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[4] ),
    .B(_02921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03659_));
 sky130_fd_sc_hd__a221o_1 _09390_ (.A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[3] ),
    .A2(_02906_),
    .B1(_03646_),
    .B2(_03647_),
    .C1(_03654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03660_));
 sky130_fd_sc_hd__or3b_2 _09391_ (.A(_03658_),
    .B(_03659_),
    .C_N(_03660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03661_));
 sky130_fd_sc_hd__a21bo_1 _09392_ (.A1(_03651_),
    .A2(_03660_),
    .B1_N(_03659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03662_));
 sky130_fd_sc_hd__a31o_1 _09393_ (.A1(_03170_),
    .A2(_03661_),
    .A3(_03662_),
    .B1(_02927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[4] ));
 sky130_fd_sc_hd__nand2_2 _09394_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[4] ),
    .B(_02921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03663_));
 sky130_fd_sc_hd__xnor2_1 _09395_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[5] ),
    .B(_02934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03664_));
 sky130_fd_sc_hd__nand3_1 _09396_ (.A(_03663_),
    .B(_03661_),
    .C(_03664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03665_));
 sky130_fd_sc_hd__a21o_1 _09397_ (.A1(_03663_),
    .A2(_03661_),
    .B1(_03664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03666_));
 sky130_fd_sc_hd__a31o_1 _09398_ (.A1(_03170_),
    .A2(_03665_),
    .A3(_03666_),
    .B1(_02943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[5] ));
 sky130_fd_sc_hd__xnor2_4 _09399_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[6] ),
    .B(_02946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03667_));
 sky130_fd_sc_hd__nand2_1 _09400_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[5] ),
    .B(_02934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03668_));
 sky130_fd_sc_hd__nor2_1 _09401_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[5] ),
    .B(_02934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03669_));
 sky130_fd_sc_hd__a31o_1 _09402_ (.A1(_03663_),
    .A2(_03661_),
    .A3(_03668_),
    .B1(_03669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03670_));
 sky130_fd_sc_hd__xor2_1 _09403_ (.A(_03667_),
    .B(_03670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03671_));
 sky130_fd_sc_hd__mux2_1 _09404_ (.A0(_02947_),
    .A1(_03671_),
    .S(_02914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03672_));
 sky130_fd_sc_hd__clkbuf_1 _09405_ (.A(_03672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[6] ));
 sky130_fd_sc_hd__a21oi_1 _09406_ (.A1(_02962_),
    .A2(_02963_),
    .B1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03673_));
 sky130_fd_sc_hd__and3_1 _09407_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[7] ),
    .B(_02962_),
    .C(_02963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03674_));
 sky130_fd_sc_hd__or2_2 _09408_ (.A(_03673_),
    .B(_03674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03675_));
 sky130_fd_sc_hd__nand2_1 _09409_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[6] ),
    .B(_02947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03676_));
 sky130_fd_sc_hd__o21ai_1 _09410_ (.A1(_03667_),
    .A2(_03670_),
    .B1(_03676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03677_));
 sky130_fd_sc_hd__xnor2_1 _09411_ (.A(_03675_),
    .B(_03677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03678_));
 sky130_fd_sc_hd__mux2_1 _09412_ (.A0(_02964_),
    .A1(_03678_),
    .S(_02853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03679_));
 sky130_fd_sc_hd__clkbuf_1 _09413_ (.A(_03679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[7] ));
 sky130_fd_sc_hd__and3_1 _09414_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[8] ),
    .B(_02975_),
    .C(_02976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03680_));
 sky130_fd_sc_hd__a21oi_1 _09415_ (.A1(_02975_),
    .A2(_02976_),
    .B1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03681_));
 sky130_fd_sc_hd__or2_1 _09416_ (.A(_03680_),
    .B(_03681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03682_));
 sky130_fd_sc_hd__and3b_1 _09417_ (.A_N(_03673_),
    .B(_02947_),
    .C(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03683_));
 sky130_fd_sc_hd__a2111oi_4 _09418_ (.A1(_03663_),
    .A2(_03668_),
    .B1(_03669_),
    .C1(_03667_),
    .D1(_03675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03684_));
 sky130_fd_sc_hd__nor4_2 _09419_ (.A(_03661_),
    .B(_03664_),
    .C(_03667_),
    .D(_03675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03685_));
 sky130_fd_sc_hd__nor4_2 _09420_ (.A(_03674_),
    .B(_03683_),
    .C(_03684_),
    .D(_03685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03686_));
 sky130_fd_sc_hd__xor2_1 _09421_ (.A(_03682_),
    .B(_03686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03687_));
 sky130_fd_sc_hd__mux2_1 _09422_ (.A0(_02978_),
    .A1(_03687_),
    .S(_02853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03688_));
 sky130_fd_sc_hd__clkbuf_1 _09423_ (.A(_03688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[8] ));
 sky130_fd_sc_hd__and3_1 _09424_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[9] ),
    .B(_02998_),
    .C(_02991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03689_));
 sky130_fd_sc_hd__a21oi_1 _09425_ (.A1(_02998_),
    .A2(_02991_),
    .B1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03690_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09426_ (.A(_03690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03691_));
 sky130_fd_sc_hd__o21ba_1 _09427_ (.A1(_03682_),
    .A2(_03686_),
    .B1_N(_03680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03692_));
 sky130_fd_sc_hd__o21ai_1 _09428_ (.A1(_03689_),
    .A2(_03691_),
    .B1(_03692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03693_));
 sky130_fd_sc_hd__o31a_1 _09429_ (.A1(_03689_),
    .A2(_03691_),
    .A3(_03692_),
    .B1(_02854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03694_));
 sky130_fd_sc_hd__a22o_1 _09430_ (.A1(_02928_),
    .A2(_02999_),
    .B1(_03693_),
    .B2(_03694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[9] ));
 sky130_fd_sc_hd__xnor2_1 _09431_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[10] ),
    .B(_03008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03695_));
 sky130_fd_sc_hd__nor2_1 _09432_ (.A(_03680_),
    .B(_03689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03696_));
 sky130_fd_sc_hd__o21a_1 _09433_ (.A1(_03682_),
    .A2(_03686_),
    .B1(_03696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03697_));
 sky130_fd_sc_hd__or3_1 _09434_ (.A(_03691_),
    .B(_03695_),
    .C(_03697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03698_));
 sky130_fd_sc_hd__o21ai_1 _09435_ (.A1(_03691_),
    .A2(_03697_),
    .B1(_03695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03699_));
 sky130_fd_sc_hd__a31o_1 _09436_ (.A1(_03170_),
    .A2(_03698_),
    .A3(_03699_),
    .B1(_03009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[10] ));
 sky130_fd_sc_hd__clkbuf_2 _09437_ (.A(_02875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03700_));
 sky130_fd_sc_hd__nand2_1 _09438_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[10] ),
    .B(_03008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03701_));
 sky130_fd_sc_hd__a21oi_1 _09439_ (.A1(_03013_),
    .A2(_03014_),
    .B1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03702_));
 sky130_fd_sc_hd__and3_1 _09440_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[11] ),
    .B(_03013_),
    .C(_03014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03703_));
 sky130_fd_sc_hd__or2_1 _09441_ (.A(_03702_),
    .B(_03703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03704_));
 sky130_fd_sc_hd__a21o_1 _09442_ (.A1(_03701_),
    .A2(_03698_),
    .B1(_03704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03705_));
 sky130_fd_sc_hd__nand3_1 _09443_ (.A(_03701_),
    .B(_03698_),
    .C(_03704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03706_));
 sky130_fd_sc_hd__a31o_1 _09444_ (.A1(_03700_),
    .A2(_03705_),
    .A3(_03706_),
    .B1(_03020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[11] ));
 sky130_fd_sc_hd__o21ba_1 _09445_ (.A1(_03701_),
    .A2(_03702_),
    .B1_N(_03703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03707_));
 sky130_fd_sc_hd__or4_1 _09446_ (.A(_03690_),
    .B(_03695_),
    .C(_03696_),
    .D(_03704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03708_));
 sky130_fd_sc_hd__or4_1 _09447_ (.A(_03680_),
    .B(_03681_),
    .C(_03689_),
    .D(_03690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03709_));
 sky130_fd_sc_hd__nor4_1 _09448_ (.A(_03695_),
    .B(_03709_),
    .C(_03702_),
    .D(_03703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03710_));
 sky130_fd_sc_hd__o41ai_2 _09449_ (.A1(_03674_),
    .A2(_03683_),
    .A3(_03684_),
    .A4(_03685_),
    .B1(_03710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03711_));
 sky130_fd_sc_hd__nand2_1 _09450_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[12] ),
    .B(_03031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03712_));
 sky130_fd_sc_hd__or2_1 _09451_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[12] ),
    .B(_03030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03713_));
 sky130_fd_sc_hd__nand2_1 _09452_ (.A(_03712_),
    .B(_03713_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03714_));
 sky130_fd_sc_hd__a31o_1 _09453_ (.A1(_03707_),
    .A2(_03708_),
    .A3(_03711_),
    .B1(_03714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03715_));
 sky130_fd_sc_hd__or4_1 _09454_ (.A(_03691_),
    .B(_03695_),
    .C(_03697_),
    .D(_03704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03716_));
 sky130_fd_sc_hd__nand3_1 _09455_ (.A(_03714_),
    .B(_03707_),
    .C(_03716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03717_));
 sky130_fd_sc_hd__a31o_1 _09456_ (.A1(_03700_),
    .A2(_03715_),
    .A3(_03717_),
    .B1(_03035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[12] ));
 sky130_fd_sc_hd__and3_1 _09457_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[13] ),
    .B(_03037_),
    .C(_03039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03718_));
 sky130_fd_sc_hd__a21oi_1 _09458_ (.A1(_03037_),
    .A2(_03039_),
    .B1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03719_));
 sky130_fd_sc_hd__nor2_1 _09459_ (.A(_03718_),
    .B(_03719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03720_));
 sky130_fd_sc_hd__and2_1 _09460_ (.A(_03712_),
    .B(_03715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03721_));
 sky130_fd_sc_hd__xnor2_1 _09461_ (.A(_03720_),
    .B(_03721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03722_));
 sky130_fd_sc_hd__a21o_1 _09462_ (.A1(_02916_),
    .A2(_03722_),
    .B1(_03045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[13] ));
 sky130_fd_sc_hd__nand2_1 _09463_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[14] ),
    .B(_03050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03723_));
 sky130_fd_sc_hd__or2_1 _09464_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[14] ),
    .B(_03050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03724_));
 sky130_fd_sc_hd__nand2_1 _09465_ (.A(_03723_),
    .B(_03724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03725_));
 sky130_fd_sc_hd__nor2_1 _09466_ (.A(_03719_),
    .B(_03721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03726_));
 sky130_fd_sc_hd__nor2_1 _09467_ (.A(_03718_),
    .B(_03726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03727_));
 sky130_fd_sc_hd__or2_1 _09468_ (.A(_03725_),
    .B(_03727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03728_));
 sky130_fd_sc_hd__a21oi_1 _09469_ (.A1(_03725_),
    .A2(_03727_),
    .B1(_02950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03729_));
 sky130_fd_sc_hd__a21o_1 _09470_ (.A1(_03728_),
    .A2(_03729_),
    .B1(_03057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[14] ));
 sky130_fd_sc_hd__and2_1 _09471_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[15] ),
    .B(_03059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03730_));
 sky130_fd_sc_hd__nor2_1 _09472_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[15] ),
    .B(_03060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03731_));
 sky130_fd_sc_hd__or2_1 _09473_ (.A(_03730_),
    .B(_03731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03732_));
 sky130_fd_sc_hd__a21o_1 _09474_ (.A1(_03723_),
    .A2(_03728_),
    .B1(_03732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03733_));
 sky130_fd_sc_hd__nand3_1 _09475_ (.A(_03723_),
    .B(_03728_),
    .C(_03732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03734_));
 sky130_fd_sc_hd__a31o_1 _09476_ (.A1(_03700_),
    .A2(_03733_),
    .A3(_03734_),
    .B1(_03066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[15] ));
 sky130_fd_sc_hd__nor2_1 _09477_ (.A(_03725_),
    .B(_03732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03735_));
 sky130_fd_sc_hd__nand2_1 _09478_ (.A(_03720_),
    .B(_03735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03736_));
 sky130_fd_sc_hd__o21bai_1 _09479_ (.A1(_03712_),
    .A2(_03719_),
    .B1_N(_03718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03737_));
 sky130_fd_sc_hd__a22oi_1 _09480_ (.A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[15] ),
    .A2(_03060_),
    .B1(_03735_),
    .B2(_03737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03738_));
 sky130_fd_sc_hd__o221a_2 _09481_ (.A1(_03723_),
    .A2(_03731_),
    .B1(_03736_),
    .B2(_03715_),
    .C1(_03738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03739_));
 sky130_fd_sc_hd__nand2_1 _09482_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[16] ),
    .B(_03117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03740_));
 sky130_fd_sc_hd__or2_1 _09483_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[16] ),
    .B(_03072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03741_));
 sky130_fd_sc_hd__nand2_1 _09484_ (.A(_03740_),
    .B(_03741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03742_));
 sky130_fd_sc_hd__or2_1 _09485_ (.A(_03739_),
    .B(_03742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03743_));
 sky130_fd_sc_hd__nand2_1 _09486_ (.A(_03739_),
    .B(_03742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03744_));
 sky130_fd_sc_hd__a31o_1 _09487_ (.A1(_03700_),
    .A2(_03743_),
    .A3(_03744_),
    .B1(_03154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[16] ));
 sky130_fd_sc_hd__o21a_1 _09488_ (.A1(_03739_),
    .A2(_03742_),
    .B1(_03740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03745_));
 sky130_fd_sc_hd__nand2_1 _09489_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[17] ),
    .B(_03098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03746_));
 sky130_fd_sc_hd__or2_1 _09490_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[17] ),
    .B(_03072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03747_));
 sky130_fd_sc_hd__nand2_1 _09491_ (.A(_03746_),
    .B(_03747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03748_));
 sky130_fd_sc_hd__xor2_1 _09492_ (.A(_03745_),
    .B(_03748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03749_));
 sky130_fd_sc_hd__clkbuf_2 _09493_ (.A(_03083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03750_));
 sky130_fd_sc_hd__a21o_1 _09494_ (.A1(_02916_),
    .A2(_03749_),
    .B1(_03750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[17] ));
 sky130_fd_sc_hd__or2b_1 _09495_ (.A(_03745_),
    .B_N(_03747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03751_));
 sky130_fd_sc_hd__nand2_1 _09496_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[18] ),
    .B(_03098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03752_));
 sky130_fd_sc_hd__or2_1 _09497_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[18] ),
    .B(_03076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03753_));
 sky130_fd_sc_hd__nand2_1 _09498_ (.A(_03752_),
    .B(_03753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03754_));
 sky130_fd_sc_hd__a21o_1 _09499_ (.A1(_03746_),
    .A2(_03751_),
    .B1(_03754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03755_));
 sky130_fd_sc_hd__nand3_1 _09500_ (.A(_03746_),
    .B(_03751_),
    .C(_03754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03756_));
 sky130_fd_sc_hd__a31o_1 _09501_ (.A1(_03700_),
    .A2(_03755_),
    .A3(_03756_),
    .B1(_03154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[18] ));
 sky130_fd_sc_hd__clkbuf_2 _09502_ (.A(_02875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03757_));
 sky130_fd_sc_hd__xnor2_1 _09503_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[19] ),
    .B(_03117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03758_));
 sky130_fd_sc_hd__a21o_1 _09504_ (.A1(_03752_),
    .A2(_03755_),
    .B1(_03758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03759_));
 sky130_fd_sc_hd__nand3_1 _09505_ (.A(_03752_),
    .B(_03755_),
    .C(_03758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03760_));
 sky130_fd_sc_hd__clkbuf_2 _09506_ (.A(_03082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03761_));
 sky130_fd_sc_hd__a31o_1 _09507_ (.A1(_03757_),
    .A2(_03759_),
    .A3(_03760_),
    .B1(_03761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[19] ));
 sky130_fd_sc_hd__o41ai_4 _09508_ (.A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[16] ),
    .A2(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[17] ),
    .A3(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[18] ),
    .A4(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[19] ),
    .B1(_03079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03762_));
 sky130_fd_sc_hd__or4_1 _09509_ (.A(_03742_),
    .B(_03748_),
    .C(_03754_),
    .D(_03758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03763_));
 sky130_fd_sc_hd__or2_1 _09510_ (.A(_03739_),
    .B(_03763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03764_));
 sky130_fd_sc_hd__nand2_1 _09511_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[20] ),
    .B(_03098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03765_));
 sky130_fd_sc_hd__or2_1 _09512_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[20] ),
    .B(_03072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03766_));
 sky130_fd_sc_hd__nand2_1 _09513_ (.A(_03765_),
    .B(_03766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03767_));
 sky130_fd_sc_hd__a21o_1 _09514_ (.A1(_03762_),
    .A2(_03764_),
    .B1(_03767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03768_));
 sky130_fd_sc_hd__a31oi_1 _09515_ (.A1(_03767_),
    .A2(_03762_),
    .A3(_03764_),
    .B1(_02950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03769_));
 sky130_fd_sc_hd__a21o_1 _09516_ (.A1(_03768_),
    .A2(_03769_),
    .B1(_03750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[20] ));
 sky130_fd_sc_hd__nand2_1 _09517_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[21] ),
    .B(_03117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03770_));
 sky130_fd_sc_hd__or2_1 _09518_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[21] ),
    .B(_03072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03771_));
 sky130_fd_sc_hd__nand2_1 _09519_ (.A(_03770_),
    .B(_03771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03772_));
 sky130_fd_sc_hd__a21oi_1 _09520_ (.A1(_03765_),
    .A2(_03768_),
    .B1(_03772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03773_));
 sky130_fd_sc_hd__a31o_1 _09521_ (.A1(_03765_),
    .A2(_03768_),
    .A3(_03772_),
    .B1(_03127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03774_));
 sky130_fd_sc_hd__o21bai_1 _09522_ (.A1(_03773_),
    .A2(_03774_),
    .B1_N(_03129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[21] ));
 sky130_fd_sc_hd__a21bo_1 _09523_ (.A1(_03765_),
    .A2(_03768_),
    .B1_N(_03771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03775_));
 sky130_fd_sc_hd__and2_1 _09524_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[22] ),
    .B(_03071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03776_));
 sky130_fd_sc_hd__nor2_1 _09525_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[22] ),
    .B(_03076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03777_));
 sky130_fd_sc_hd__or2_1 _09526_ (.A(_03776_),
    .B(_03777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03778_));
 sky130_fd_sc_hd__a21oi_1 _09527_ (.A1(_03770_),
    .A2(_03775_),
    .B1(_03778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03779_));
 sky130_fd_sc_hd__a31o_1 _09528_ (.A1(_03770_),
    .A2(_03775_),
    .A3(_03778_),
    .B1(_03127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03780_));
 sky130_fd_sc_hd__o21bai_1 _09529_ (.A1(_03779_),
    .A2(_03780_),
    .B1_N(_03129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[22] ));
 sky130_fd_sc_hd__xor2_1 _09530_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[23] ),
    .B(_03117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03781_));
 sky130_fd_sc_hd__o21ai_1 _09531_ (.A1(_03776_),
    .A2(_03779_),
    .B1(_03781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03782_));
 sky130_fd_sc_hd__or3_1 _09532_ (.A(_03776_),
    .B(_03779_),
    .C(_03781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03783_));
 sky130_fd_sc_hd__a31o_1 _09533_ (.A1(_03757_),
    .A2(_03782_),
    .A3(_03783_),
    .B1(_03761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[23] ));
 sky130_fd_sc_hd__or4b_1 _09534_ (.A(_03767_),
    .B(_03772_),
    .C(_03778_),
    .D_N(_03781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03784_));
 sky130_fd_sc_hd__or2_1 _09535_ (.A(_03763_),
    .B(_03784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03785_));
 sky130_fd_sc_hd__o41ai_4 _09536_ (.A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[20] ),
    .A2(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[21] ),
    .A3(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[22] ),
    .A4(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[23] ),
    .B1(_03079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03786_));
 sky130_fd_sc_hd__o211ai_4 _09537_ (.A1(_03739_),
    .A2(_03785_),
    .B1(_03786_),
    .C1(_03762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03787_));
 sky130_fd_sc_hd__xor2_1 _09538_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[24] ),
    .B(_03138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03788_));
 sky130_fd_sc_hd__nand2_1 _09539_ (.A(_03787_),
    .B(_03788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03789_));
 sky130_fd_sc_hd__o21a_1 _09540_ (.A1(_03787_),
    .A2(_03788_),
    .B1(_02877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03790_));
 sky130_fd_sc_hd__a21o_1 _09541_ (.A1(_03789_),
    .A2(_03790_),
    .B1(_03750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[24] ));
 sky130_fd_sc_hd__xor2_1 _09542_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[25] ),
    .B(_03138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03791_));
 sky130_fd_sc_hd__a22o_1 _09543_ (.A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[24] ),
    .A2(_03143_),
    .B1(_03787_),
    .B2(_03788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03792_));
 sky130_fd_sc_hd__xor2_1 _09544_ (.A(_03791_),
    .B(_03792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03793_));
 sky130_fd_sc_hd__a21o_1 _09545_ (.A1(_02916_),
    .A2(_03793_),
    .B1(_03750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[25] ));
 sky130_fd_sc_hd__o21ai_1 _09546_ (.A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[24] ),
    .A2(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[25] ),
    .B1(_03081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03794_));
 sky130_fd_sc_hd__and2_1 _09547_ (.A(_03788_),
    .B(_03791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03795_));
 sky130_fd_sc_hd__nand2_1 _09548_ (.A(_03787_),
    .B(_03795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03796_));
 sky130_fd_sc_hd__nand2_1 _09549_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[26] ),
    .B(_03085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03797_));
 sky130_fd_sc_hd__or2_1 _09550_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[26] ),
    .B(_03078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03798_));
 sky130_fd_sc_hd__nand2_1 _09551_ (.A(_03797_),
    .B(_03798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03799_));
 sky130_fd_sc_hd__a21o_1 _09552_ (.A1(_03794_),
    .A2(_03796_),
    .B1(_03799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03800_));
 sky130_fd_sc_hd__nand3_1 _09553_ (.A(_03799_),
    .B(_03794_),
    .C(_03796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03801_));
 sky130_fd_sc_hd__a31o_1 _09554_ (.A1(_03757_),
    .A2(_03800_),
    .A3(_03801_),
    .B1(_03761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[26] ));
 sky130_fd_sc_hd__xnor2_1 _09555_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[27] ),
    .B(_03085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03802_));
 sky130_fd_sc_hd__nand2_1 _09556_ (.A(_03797_),
    .B(_03800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03803_));
 sky130_fd_sc_hd__xnor2_1 _09557_ (.A(_03802_),
    .B(_03803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03804_));
 sky130_fd_sc_hd__a21o_1 _09558_ (.A1(_02916_),
    .A2(_03804_),
    .B1(_03750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[27] ));
 sky130_fd_sc_hd__nor2_1 _09559_ (.A(_03799_),
    .B(_03802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03805_));
 sky130_fd_sc_hd__o41a_1 _09560_ (.A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[24] ),
    .A2(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[25] ),
    .A3(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[26] ),
    .A4(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[27] ),
    .B1(_03086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03806_));
 sky130_fd_sc_hd__a31oi_2 _09561_ (.A1(_03787_),
    .A2(_03795_),
    .A3(_03805_),
    .B1(_03806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03807_));
 sky130_fd_sc_hd__and2_1 _09562_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[28] ),
    .B(_03079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03808_));
 sky130_fd_sc_hd__nor2_1 _09563_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[28] ),
    .B(_03086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03809_));
 sky130_fd_sc_hd__or2_1 _09564_ (.A(_03808_),
    .B(_03809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03810_));
 sky130_fd_sc_hd__nor2_1 _09565_ (.A(_03807_),
    .B(_03810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03811_));
 sky130_fd_sc_hd__a21o_1 _09566_ (.A1(_03807_),
    .A2(_03810_),
    .B1(_03127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03812_));
 sky130_fd_sc_hd__o21bai_1 _09567_ (.A1(_03811_),
    .A2(_03812_),
    .B1_N(_03083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[28] ));
 sky130_fd_sc_hd__nand2_1 _09568_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[29] ),
    .B(_03080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03813_));
 sky130_fd_sc_hd__or2_1 _09569_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[29] ),
    .B(_03080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03814_));
 sky130_fd_sc_hd__o211ai_1 _09570_ (.A1(_03808_),
    .A2(_03811_),
    .B1(_03813_),
    .C1(_03814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03815_));
 sky130_fd_sc_hd__a211o_1 _09571_ (.A1(_03813_),
    .A2(_03814_),
    .B1(_03808_),
    .C1(_03811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03816_));
 sky130_fd_sc_hd__a31o_1 _09572_ (.A1(_03757_),
    .A2(_03815_),
    .A3(_03816_),
    .B1(_03761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[29] ));
 sky130_fd_sc_hd__o21ai_1 _09573_ (.A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[28] ),
    .A2(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[29] ),
    .B1(_03081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03817_));
 sky130_fd_sc_hd__or4bb_1 _09574_ (.A(_03807_),
    .B(_03810_),
    .C_N(_03813_),
    .D_N(_03814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03818_));
 sky130_fd_sc_hd__nand2_1 _09575_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[30] ),
    .B(_03087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03819_));
 sky130_fd_sc_hd__or2_1 _09576_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[30] ),
    .B(_03087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03820_));
 sky130_fd_sc_hd__nand2_1 _09577_ (.A(_03819_),
    .B(_03820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03821_));
 sky130_fd_sc_hd__a21o_1 _09578_ (.A1(_03817_),
    .A2(_03818_),
    .B1(_03821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03822_));
 sky130_fd_sc_hd__nand3_1 _09579_ (.A(_03821_),
    .B(_03817_),
    .C(_03818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03823_));
 sky130_fd_sc_hd__a31o_1 _09580_ (.A1(_03757_),
    .A2(_03822_),
    .A3(_03823_),
    .B1(_03761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[30] ));
 sky130_fd_sc_hd__xnor2_1 _09581_ (.A(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[31] ),
    .B(_03143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03824_));
 sky130_fd_sc_hd__a21oi_1 _09582_ (.A1(_03819_),
    .A2(_03822_),
    .B1(_03824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03825_));
 sky130_fd_sc_hd__a31o_1 _09583_ (.A1(_03819_),
    .A2(_03822_),
    .A3(_03824_),
    .B1(_02898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03826_));
 sky130_fd_sc_hd__o21bai_1 _09584_ (.A1(_03825_),
    .A2(_03826_),
    .B1_N(_03083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[31] ));
 sky130_fd_sc_hd__mux2_1 _09585_ (.A0(\sa_inst.sak._17_[0] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[0] ),
    .S(_03419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03827_));
 sky130_fd_sc_hd__clkbuf_2 _09586_ (.A(_03827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ));
 sky130_fd_sc_hd__mux2_1 _09587_ (.A0(\sa_inst.sak._17_[1] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[1] ),
    .S(_03419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03828_));
 sky130_fd_sc_hd__buf_2 _09588_ (.A(_03828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ));
 sky130_fd_sc_hd__clkbuf_2 _09589_ (.A(_03406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03829_));
 sky130_fd_sc_hd__mux2_1 _09590_ (.A0(\sa_inst.sak._17_[2] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[2] ),
    .S(_03829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03830_));
 sky130_fd_sc_hd__clkbuf_2 _09591_ (.A(_03830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ));
 sky130_fd_sc_hd__mux2_2 _09592_ (.A0(\sa_inst.sak._17_[3] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[3] ),
    .S(_03829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03831_));
 sky130_fd_sc_hd__clkbuf_1 _09593_ (.A(_03831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ));
 sky130_fd_sc_hd__mux2_1 _09594_ (.A0(\sa_inst.sak._17_[4] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[4] ),
    .S(_03829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03832_));
 sky130_fd_sc_hd__clkbuf_2 _09595_ (.A(_03832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ));
 sky130_fd_sc_hd__mux2_2 _09596_ (.A0(\sa_inst.sak._17_[5] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[5] ),
    .S(_03829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03833_));
 sky130_fd_sc_hd__clkbuf_1 _09597_ (.A(_03833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ));
 sky130_fd_sc_hd__mux2_2 _09598_ (.A0(\sa_inst.sak._17_[6] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[6] ),
    .S(_03829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03834_));
 sky130_fd_sc_hd__clkbuf_1 _09599_ (.A(_03834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ));
 sky130_fd_sc_hd__clkbuf_2 _09600_ (.A(_03406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03835_));
 sky130_fd_sc_hd__mux2_2 _09601_ (.A0(\sa_inst.sak._17_[7] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[7] ),
    .S(_03835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03836_));
 sky130_fd_sc_hd__clkbuf_1 _09602_ (.A(_03836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ));
 sky130_fd_sc_hd__mux2_2 _09603_ (.A0(\sa_inst.sak._17_[8] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[8] ),
    .S(_03835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03837_));
 sky130_fd_sc_hd__clkbuf_1 _09604_ (.A(_03837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ));
 sky130_fd_sc_hd__mux2_2 _09605_ (.A0(\sa_inst.sak._17_[9] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[9] ),
    .S(_03835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03838_));
 sky130_fd_sc_hd__clkbuf_1 _09606_ (.A(_03838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ));
 sky130_fd_sc_hd__mux2_2 _09607_ (.A0(\sa_inst.sak._17_[10] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[10] ),
    .S(_03835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03839_));
 sky130_fd_sc_hd__clkbuf_1 _09608_ (.A(_03839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ));
 sky130_fd_sc_hd__mux2_2 _09609_ (.A0(\sa_inst.sak._17_[11] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[11] ),
    .S(_03835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03840_));
 sky130_fd_sc_hd__clkbuf_1 _09610_ (.A(_03840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ));
 sky130_fd_sc_hd__clkbuf_2 _09611_ (.A(_03405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03841_));
 sky130_fd_sc_hd__mux2_2 _09612_ (.A0(\sa_inst.sak._17_[12] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[12] ),
    .S(_03841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03842_));
 sky130_fd_sc_hd__clkbuf_1 _09613_ (.A(_03842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ));
 sky130_fd_sc_hd__mux2_1 _09614_ (.A0(\sa_inst.sak._17_[13] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[13] ),
    .S(_03841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03843_));
 sky130_fd_sc_hd__clkbuf_1 _09615_ (.A(_03843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ));
 sky130_fd_sc_hd__mux2_1 _09616_ (.A0(\sa_inst.sak._17_[14] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[14] ),
    .S(_03841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03844_));
 sky130_fd_sc_hd__clkbuf_1 _09617_ (.A(_03844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ));
 sky130_fd_sc_hd__mux2_1 _09618_ (.A0(\sa_inst.sak._17_[15] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[15] ),
    .S(_03841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03845_));
 sky130_fd_sc_hd__clkbuf_1 _09619_ (.A(_03845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ));
 sky130_fd_sc_hd__mux2_1 _09620_ (.A0(\sa_inst.sak._17_[16] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[16] ),
    .S(_03841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03846_));
 sky130_fd_sc_hd__clkbuf_1 _09621_ (.A(_03846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ));
 sky130_fd_sc_hd__clkbuf_2 _09622_ (.A(_03405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03847_));
 sky130_fd_sc_hd__mux2_1 _09623_ (.A0(\sa_inst.sak._17_[17] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[17] ),
    .S(_03847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03848_));
 sky130_fd_sc_hd__clkbuf_1 _09624_ (.A(_03848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ));
 sky130_fd_sc_hd__mux2_1 _09625_ (.A0(\sa_inst.sak._17_[18] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[18] ),
    .S(_03847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03849_));
 sky130_fd_sc_hd__clkbuf_1 _09626_ (.A(_03849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ));
 sky130_fd_sc_hd__mux2_1 _09627_ (.A0(\sa_inst.sak._17_[19] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[19] ),
    .S(_03847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03850_));
 sky130_fd_sc_hd__clkbuf_1 _09628_ (.A(_03850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ));
 sky130_fd_sc_hd__mux2_1 _09629_ (.A0(\sa_inst.sak._17_[20] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[20] ),
    .S(_03847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03851_));
 sky130_fd_sc_hd__clkbuf_1 _09630_ (.A(_03851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ));
 sky130_fd_sc_hd__mux2_1 _09631_ (.A0(\sa_inst.sak._17_[21] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[21] ),
    .S(_03847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03852_));
 sky130_fd_sc_hd__clkbuf_1 _09632_ (.A(_03852_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ));
 sky130_fd_sc_hd__clkbuf_2 _09633_ (.A(_03405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03853_));
 sky130_fd_sc_hd__mux2_1 _09634_ (.A0(\sa_inst.sak._17_[22] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[22] ),
    .S(_03853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03854_));
 sky130_fd_sc_hd__clkbuf_1 _09635_ (.A(_03854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ));
 sky130_fd_sc_hd__mux2_1 _09636_ (.A0(\sa_inst.sak._17_[23] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[23] ),
    .S(_03853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03855_));
 sky130_fd_sc_hd__clkbuf_1 _09637_ (.A(_03855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ));
 sky130_fd_sc_hd__mux2_1 _09638_ (.A0(\sa_inst.sak._17_[24] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[24] ),
    .S(_03853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03856_));
 sky130_fd_sc_hd__clkbuf_1 _09639_ (.A(_03856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ));
 sky130_fd_sc_hd__mux2_1 _09640_ (.A0(\sa_inst.sak._17_[25] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[25] ),
    .S(_03853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03857_));
 sky130_fd_sc_hd__clkbuf_1 _09641_ (.A(_03857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ));
 sky130_fd_sc_hd__mux2_1 _09642_ (.A0(\sa_inst.sak._17_[26] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[26] ),
    .S(_03853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03858_));
 sky130_fd_sc_hd__clkbuf_1 _09643_ (.A(_03858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ));
 sky130_fd_sc_hd__clkbuf_2 _09644_ (.A(_03405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03859_));
 sky130_fd_sc_hd__mux2_1 _09645_ (.A0(\sa_inst.sak._17_[27] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[27] ),
    .S(_03859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03860_));
 sky130_fd_sc_hd__clkbuf_1 _09646_ (.A(_03860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ));
 sky130_fd_sc_hd__mux2_1 _09647_ (.A0(\sa_inst.sak._17_[28] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[28] ),
    .S(_03859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03861_));
 sky130_fd_sc_hd__clkbuf_1 _09648_ (.A(_03861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ));
 sky130_fd_sc_hd__mux2_1 _09649_ (.A0(\sa_inst.sak._17_[29] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[29] ),
    .S(_03859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03862_));
 sky130_fd_sc_hd__clkbuf_1 _09650_ (.A(_03862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ));
 sky130_fd_sc_hd__mux2_1 _09651_ (.A0(\sa_inst.sak._17_[30] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[30] ),
    .S(_03859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03863_));
 sky130_fd_sc_hd__clkbuf_1 _09652_ (.A(_03863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ));
 sky130_fd_sc_hd__mux2_1 _09653_ (.A0(\sa_inst.sak._17_[31] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[31] ),
    .S(_03859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03864_));
 sky130_fd_sc_hd__clkbuf_1 _09654_ (.A(_03864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ));
 sky130_fd_sc_hd__mux2_1 _09655_ (.A0(\sa_inst.sak._17_[32] ),
    .A1(\sa_inst.sak.rows:3.cols:2.pe_ij._02_ ),
    .S(_03380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03865_));
 sky130_fd_sc_hd__buf_2 _09656_ (.A(_03865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ));
 sky130_fd_sc_hd__inv_2 _09657_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._22_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03866_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09658_ (.A(_03866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03867_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09659_ (.A(_03867_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03868_));
 sky130_fd_sc_hd__inv_2 _09660_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03869_));
 sky130_fd_sc_hd__clkbuf_2 _09661_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03870_));
 sky130_fd_sc_hd__mux4_2 _09662_ (.A0(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .A2(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .A3(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .S0(_03870_),
    .S1(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03871_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09663_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03872_));
 sky130_fd_sc_hd__mux2_1 _09664_ (.A0(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[1] ),
    .S(_03872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03873_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09665_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03874_));
 sky130_fd_sc_hd__and2b_1 _09666_ (.A_N(_03874_),
    .B(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03875_));
 sky130_fd_sc_hd__a22o_1 _09667_ (.A1(_03869_),
    .A2(_03871_),
    .B1(_03873_),
    .B2(_03875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03876_));
 sky130_fd_sc_hd__nand2_1 _09668_ (.A(_03868_),
    .B(_03876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03877_));
 sky130_fd_sc_hd__buf_4 _09669_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03878_));
 sky130_fd_sc_hd__nand2_1 _09670_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[0] ),
    .B(_03878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03879_));
 sky130_fd_sc_hd__xor2_1 _09671_ (.A(_03877_),
    .B(_03879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[0] ));
 sky130_fd_sc_hd__inv_2 _09672_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03880_));
 sky130_fd_sc_hd__or2b_1 _09673_ (.A(_03874_),
    .B_N(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03881_));
 sky130_fd_sc_hd__clkbuf_2 _09674_ (.A(_03870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03882_));
 sky130_fd_sc_hd__or2b_1 _09675_ (.A(_03882_),
    .B_N(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03883_));
 sky130_fd_sc_hd__mux4_2 _09676_ (.A0(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .A2(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .A3(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .S0(_03870_),
    .S1(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03884_));
 sky130_fd_sc_hd__a2bb2o_1 _09677_ (.A1_N(_03881_),
    .A2_N(_03883_),
    .B1(_03884_),
    .B2(_03869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03885_));
 sky130_fd_sc_hd__and3_1 _09678_ (.A(_03866_),
    .B(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[0] ),
    .C(_03876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03886_));
 sky130_fd_sc_hd__and3_1 _09679_ (.A(_03866_),
    .B(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[1] ),
    .C(_03885_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03887_));
 sky130_fd_sc_hd__a21o_1 _09680_ (.A1(_03867_),
    .A2(_03885_),
    .B1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03888_));
 sky130_fd_sc_hd__or2b_1 _09681_ (.A(_03887_),
    .B_N(_03888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03889_));
 sky130_fd_sc_hd__xnor2_1 _09682_ (.A(_03886_),
    .B(_03889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03890_));
 sky130_fd_sc_hd__and2_1 _09683_ (.A(_03878_),
    .B(_03890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03891_));
 sky130_fd_sc_hd__a31o_1 _09684_ (.A1(_03868_),
    .A2(_03880_),
    .A3(_03885_),
    .B1(_03891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[1] ));
 sky130_fd_sc_hd__mux2_1 _09685_ (.A0(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .S(_03870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03892_));
 sky130_fd_sc_hd__and2_1 _09686_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .B(_03872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03893_));
 sky130_fd_sc_hd__and2b_1 _09687_ (.A_N(_03872_),
    .B(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03894_));
 sky130_fd_sc_hd__mux2_1 _09688_ (.A0(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ),
    .S(_03870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03895_));
 sky130_fd_sc_hd__inv_2 _09689_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03896_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09690_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03897_));
 sky130_fd_sc_hd__mux4_1 _09691_ (.A0(_03892_),
    .A1(_03893_),
    .A2(_03894_),
    .A3(_03895_),
    .S0(_03896_),
    .S1(_03897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03898_));
 sky130_fd_sc_hd__and2_1 _09692_ (.A(_03866_),
    .B(_03898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03899_));
 sky130_fd_sc_hd__a21o_1 _09693_ (.A1(_03886_),
    .A2(_03888_),
    .B1(_03887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03900_));
 sky130_fd_sc_hd__or2_1 _09694_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[2] ),
    .B(_03899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03901_));
 sky130_fd_sc_hd__nand2_1 _09695_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[2] ),
    .B(_03899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03902_));
 sky130_fd_sc_hd__nand2_1 _09696_ (.A(_03901_),
    .B(_03902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03903_));
 sky130_fd_sc_hd__xnor2_1 _09697_ (.A(_03900_),
    .B(_03903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03904_));
 sky130_fd_sc_hd__mux2_1 _09698_ (.A0(_03899_),
    .A1(_03904_),
    .S(_03878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03905_));
 sky130_fd_sc_hd__clkbuf_1 _09699_ (.A(_03905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[2] ));
 sky130_fd_sc_hd__mux2_1 _09700_ (.A0(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .S(_03882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03906_));
 sky130_fd_sc_hd__a21o_1 _09701_ (.A1(_03882_),
    .A2(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .B1(_03874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03907_));
 sky130_fd_sc_hd__o211a_1 _09702_ (.A1(_03896_),
    .A2(_03906_),
    .B1(_03907_),
    .C1(_03869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03908_));
 sky130_fd_sc_hd__mux2_1 _09703_ (.A0(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ),
    .S(_03882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03909_));
 sky130_fd_sc_hd__and2_1 _09704_ (.A(_03875_),
    .B(_03909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03910_));
 sky130_fd_sc_hd__o21a_1 _09705_ (.A1(_03908_),
    .A2(_03910_),
    .B1(_03867_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03911_));
 sky130_fd_sc_hd__nor2_1 _09706_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[3] ),
    .B(_03911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03912_));
 sky130_fd_sc_hd__and2_1 _09707_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[3] ),
    .B(_03911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03913_));
 sky130_fd_sc_hd__or2_1 _09708_ (.A(_03912_),
    .B(_03913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03914_));
 sky130_fd_sc_hd__and3_1 _09709_ (.A(_03868_),
    .B(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[2] ),
    .C(_03898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03915_));
 sky130_fd_sc_hd__a21o_1 _09710_ (.A1(_03900_),
    .A2(_03901_),
    .B1(_03915_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03916_));
 sky130_fd_sc_hd__xnor2_1 _09711_ (.A(_03914_),
    .B(_03916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03917_));
 sky130_fd_sc_hd__mux2_1 _09712_ (.A0(_03911_),
    .A1(_03917_),
    .S(_03878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03918_));
 sky130_fd_sc_hd__clkbuf_1 _09713_ (.A(_03918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[3] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09714_ (.A(_03874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03919_));
 sky130_fd_sc_hd__mux2_1 _09715_ (.A0(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ),
    .S(_03882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03920_));
 sky130_fd_sc_hd__a21o_1 _09716_ (.A1(_03919_),
    .A2(_03920_),
    .B1(_03897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03921_));
 sky130_fd_sc_hd__mux2_1 _09717_ (.A0(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ),
    .S(_03872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03922_));
 sky130_fd_sc_hd__nand2_1 _09718_ (.A(_03874_),
    .B(_03897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03923_));
 sky130_fd_sc_hd__o22a_1 _09719_ (.A1(_03922_),
    .A2(_03881_),
    .B1(_03923_),
    .B2(_03873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03924_));
 sky130_fd_sc_hd__and3_1 _09720_ (.A(_03866_),
    .B(_03921_),
    .C(_03924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03925_));
 sky130_fd_sc_hd__nand2_1 _09721_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[4] ),
    .B(_03925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03926_));
 sky130_fd_sc_hd__or2_1 _09722_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[4] ),
    .B(_03925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03927_));
 sky130_fd_sc_hd__nand2_1 _09723_ (.A(_03926_),
    .B(_03927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03928_));
 sky130_fd_sc_hd__a211oi_1 _09724_ (.A1(_03900_),
    .A2(_03901_),
    .B1(_03915_),
    .C1(_03913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03929_));
 sky130_fd_sc_hd__or2_1 _09725_ (.A(_03912_),
    .B(_03929_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03930_));
 sky130_fd_sc_hd__xor2_1 _09726_ (.A(_03928_),
    .B(_03930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03931_));
 sky130_fd_sc_hd__clkbuf_2 _09727_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03932_));
 sky130_fd_sc_hd__buf_2 _09728_ (.A(_03932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03933_));
 sky130_fd_sc_hd__mux2_1 _09729_ (.A0(_03925_),
    .A1(_03931_),
    .S(_03933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03934_));
 sky130_fd_sc_hd__clkbuf_1 _09730_ (.A(_03934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[4] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09731_ (.A(_03872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03935_));
 sky130_fd_sc_hd__mux2_1 _09732_ (.A0(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ),
    .S(_03935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03936_));
 sky130_fd_sc_hd__mux2_1 _09733_ (.A0(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ),
    .S(_03935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03937_));
 sky130_fd_sc_hd__a21o_1 _09734_ (.A1(_03919_),
    .A2(_03937_),
    .B1(_03897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03938_));
 sky130_fd_sc_hd__clkbuf_1 _09735_ (.A(_03919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03939_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09736_ (.A(_03897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03940_));
 sky130_fd_sc_hd__a31oi_1 _09737_ (.A1(_03939_),
    .A2(_03940_),
    .A3(_03883_),
    .B1(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._22_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03941_));
 sky130_fd_sc_hd__o211a_1 _09738_ (.A1(_03881_),
    .A2(_03936_),
    .B1(_03938_),
    .C1(_03941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03942_));
 sky130_fd_sc_hd__xnor2_1 _09739_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[5] ),
    .B(_03942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03943_));
 sky130_fd_sc_hd__o21a_1 _09740_ (.A1(_03928_),
    .A2(_03930_),
    .B1(_03926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03944_));
 sky130_fd_sc_hd__xor2_1 _09741_ (.A(_03943_),
    .B(_03944_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03945_));
 sky130_fd_sc_hd__mux2_1 _09742_ (.A0(_03942_),
    .A1(_03945_),
    .S(_03933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03946_));
 sky130_fd_sc_hd__clkbuf_1 _09743_ (.A(_03946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[5] ));
 sky130_fd_sc_hd__o22a_1 _09744_ (.A1(_03881_),
    .A2(_03892_),
    .B1(_03895_),
    .B2(_03923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03947_));
 sky130_fd_sc_hd__a31o_1 _09745_ (.A1(_03919_),
    .A2(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ),
    .A3(_03935_),
    .B1(_03940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03948_));
 sky130_fd_sc_hd__and3_1 _09746_ (.A(_03867_),
    .B(_03947_),
    .C(_03948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03949_));
 sky130_fd_sc_hd__and2_1 _09747_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[6] ),
    .B(_03949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03950_));
 sky130_fd_sc_hd__nor2_1 _09748_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[6] ),
    .B(_03949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03951_));
 sky130_fd_sc_hd__or2_2 _09749_ (.A(_03950_),
    .B(_03951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03952_));
 sky130_fd_sc_hd__a22o_1 _09750_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[4] ),
    .A2(_03925_),
    .B1(_03942_),
    .B2(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03953_));
 sky130_fd_sc_hd__o21ai_1 _09751_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[5] ),
    .A2(_03942_),
    .B1(_03953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03954_));
 sky130_fd_sc_hd__o41a_2 _09752_ (.A1(_03912_),
    .A2(_03928_),
    .A3(_03929_),
    .A4(_03943_),
    .B1(_03954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03955_));
 sky130_fd_sc_hd__xor2_1 _09753_ (.A(_03952_),
    .B(_03955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03956_));
 sky130_fd_sc_hd__mux2_1 _09754_ (.A0(_03949_),
    .A1(_03956_),
    .S(_03933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03957_));
 sky130_fd_sc_hd__clkbuf_1 _09755_ (.A(_03957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[6] ));
 sky130_fd_sc_hd__o22a_1 _09756_ (.A1(_03881_),
    .A2(_03906_),
    .B1(_03909_),
    .B2(_03923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03958_));
 sky130_fd_sc_hd__a31o_1 _09757_ (.A1(_03919_),
    .A2(_03935_),
    .A3(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .B1(_03940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03959_));
 sky130_fd_sc_hd__and3_1 _09758_ (.A(_03867_),
    .B(_03958_),
    .C(_03959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03960_));
 sky130_fd_sc_hd__and2_1 _09759_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[7] ),
    .B(_03960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03961_));
 sky130_fd_sc_hd__nor2_1 _09760_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[7] ),
    .B(_03960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03962_));
 sky130_fd_sc_hd__or2_1 _09761_ (.A(_03961_),
    .B(_03962_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03963_));
 sky130_fd_sc_hd__o21bai_1 _09762_ (.A1(_03952_),
    .A2(_03955_),
    .B1_N(_03950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03964_));
 sky130_fd_sc_hd__xnor2_1 _09763_ (.A(_03963_),
    .B(_03964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03965_));
 sky130_fd_sc_hd__mux2_1 _09764_ (.A0(_03960_),
    .A1(_03965_),
    .S(_03933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03966_));
 sky130_fd_sc_hd__clkbuf_1 _09765_ (.A(_03966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[7] ));
 sky130_fd_sc_hd__and3_1 _09766_ (.A(_03940_),
    .B(_03868_),
    .C(_03871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03967_));
 sky130_fd_sc_hd__nor2_2 _09767_ (.A(_03869_),
    .B(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._22_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03968_));
 sky130_fd_sc_hd__and3_1 _09768_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[8] ),
    .B(_03871_),
    .C(_03968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03969_));
 sky130_fd_sc_hd__nor2_1 _09769_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[8] ),
    .B(_03967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03970_));
 sky130_fd_sc_hd__or2_1 _09770_ (.A(_03969_),
    .B(_03970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03971_));
 sky130_fd_sc_hd__o21bai_1 _09771_ (.A1(_03950_),
    .A2(_03961_),
    .B1_N(_03962_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03972_));
 sky130_fd_sc_hd__o31ai_4 _09772_ (.A1(_03952_),
    .A2(_03955_),
    .A3(_03963_),
    .B1(_03972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03973_));
 sky130_fd_sc_hd__xnor2_1 _09773_ (.A(_03971_),
    .B(_03973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03974_));
 sky130_fd_sc_hd__mux2_1 _09774_ (.A0(_03967_),
    .A1(_03974_),
    .S(_03933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03975_));
 sky130_fd_sc_hd__clkbuf_1 _09775_ (.A(_03975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[8] ));
 sky130_fd_sc_hd__buf_2 _09776_ (.A(_03932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03976_));
 sky130_fd_sc_hd__and3_1 _09777_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[9] ),
    .B(_03884_),
    .C(_03968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03977_));
 sky130_fd_sc_hd__and3_1 _09778_ (.A(_03940_),
    .B(_03868_),
    .C(_03884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03978_));
 sky130_fd_sc_hd__nor2_1 _09779_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[9] ),
    .B(_03978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03979_));
 sky130_fd_sc_hd__or2_1 _09780_ (.A(_03977_),
    .B(_03979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03980_));
 sky130_fd_sc_hd__inv_2 _09781_ (.A(_03971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03981_));
 sky130_fd_sc_hd__a21oi_1 _09782_ (.A1(_03981_),
    .A2(_03973_),
    .B1(_03969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03982_));
 sky130_fd_sc_hd__xnor2_1 _09783_ (.A(_03980_),
    .B(_03982_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03983_));
 sky130_fd_sc_hd__buf_2 _09784_ (.A(_03932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03984_));
 sky130_fd_sc_hd__nor2_1 _09785_ (.A(_03984_),
    .B(_03978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03985_));
 sky130_fd_sc_hd__a21oi_1 _09786_ (.A1(_03976_),
    .A2(_03983_),
    .B1(_03985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[9] ));
 sky130_fd_sc_hd__mux2_1 _09787_ (.A0(_03892_),
    .A1(_03893_),
    .S(_03896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03986_));
 sky130_fd_sc_hd__and2_1 _09788_ (.A(_03986_),
    .B(_03968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03987_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09789_ (.A(_03968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03988_));
 sky130_fd_sc_hd__and3_1 _09790_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[10] ),
    .B(_03986_),
    .C(_03988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03989_));
 sky130_fd_sc_hd__nor2_1 _09791_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[10] ),
    .B(_03987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03990_));
 sky130_fd_sc_hd__or2_1 _09792_ (.A(_03989_),
    .B(_03990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03991_));
 sky130_fd_sc_hd__inv_2 _09793_ (.A(_03979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03992_));
 sky130_fd_sc_hd__a211o_1 _09794_ (.A1(_03981_),
    .A2(_03973_),
    .B1(_03977_),
    .C1(_03969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03993_));
 sky130_fd_sc_hd__and2_1 _09795_ (.A(_03992_),
    .B(_03993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03994_));
 sky130_fd_sc_hd__xnor2_1 _09796_ (.A(_03991_),
    .B(_03994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03995_));
 sky130_fd_sc_hd__clkbuf_2 _09797_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03996_));
 sky130_fd_sc_hd__mux2_1 _09798_ (.A0(_03987_),
    .A1(_03995_),
    .S(_03996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03997_));
 sky130_fd_sc_hd__clkbuf_1 _09799_ (.A(_03997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[10] ));
 sky130_fd_sc_hd__o211a_1 _09800_ (.A1(_03896_),
    .A2(_03906_),
    .B1(_03907_),
    .C1(_03988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03998_));
 sky130_fd_sc_hd__and2_1 _09801_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[11] ),
    .B(_03998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03999_));
 sky130_fd_sc_hd__or2_1 _09802_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[11] ),
    .B(_03998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04000_));
 sky130_fd_sc_hd__or2b_1 _09803_ (.A(_03999_),
    .B_N(_04000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04001_));
 sky130_fd_sc_hd__inv_2 _09804_ (.A(_03990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04002_));
 sky130_fd_sc_hd__a31o_1 _09805_ (.A1(_03992_),
    .A2(_04002_),
    .A3(_03993_),
    .B1(_03989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04003_));
 sky130_fd_sc_hd__xnor2_1 _09806_ (.A(_04001_),
    .B(_04003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04004_));
 sky130_fd_sc_hd__mux2_1 _09807_ (.A0(_03998_),
    .A1(_04004_),
    .S(_03996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04005_));
 sky130_fd_sc_hd__clkbuf_1 _09808_ (.A(_04005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[11] ));
 sky130_fd_sc_hd__and3_1 _09809_ (.A(_03939_),
    .B(_03920_),
    .C(_03968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04006_));
 sky130_fd_sc_hd__and2_1 _09810_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[12] ),
    .B(_04006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04007_));
 sky130_fd_sc_hd__nor2_1 _09811_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[12] ),
    .B(_04006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04008_));
 sky130_fd_sc_hd__or2_1 _09812_ (.A(_04007_),
    .B(_04008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04009_));
 sky130_fd_sc_hd__inv_2 _09813_ (.A(_04009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04010_));
 sky130_fd_sc_hd__a311o_1 _09814_ (.A1(_03992_),
    .A2(_04002_),
    .A3(_03993_),
    .B1(_03999_),
    .C1(_03989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04011_));
 sky130_fd_sc_hd__nand2_1 _09815_ (.A(_04000_),
    .B(_04011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04012_));
 sky130_fd_sc_hd__xnor2_1 _09816_ (.A(_04010_),
    .B(_04012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04013_));
 sky130_fd_sc_hd__mux2_1 _09817_ (.A0(_04006_),
    .A1(_04013_),
    .S(_03996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04014_));
 sky130_fd_sc_hd__clkbuf_1 _09818_ (.A(_04014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[12] ));
 sky130_fd_sc_hd__and3_1 _09819_ (.A(_03939_),
    .B(_03937_),
    .C(_03988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04015_));
 sky130_fd_sc_hd__and2_1 _09820_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[13] ),
    .B(_04015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04016_));
 sky130_fd_sc_hd__nor2_1 _09821_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[13] ),
    .B(_04015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04017_));
 sky130_fd_sc_hd__nor2_1 _09822_ (.A(_04016_),
    .B(_04017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04018_));
 sky130_fd_sc_hd__a31o_1 _09823_ (.A1(_04000_),
    .A2(_04010_),
    .A3(_04011_),
    .B1(_04007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04019_));
 sky130_fd_sc_hd__xor2_1 _09824_ (.A(_04018_),
    .B(_04019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04020_));
 sky130_fd_sc_hd__mux2_1 _09825_ (.A0(_04015_),
    .A1(_04020_),
    .S(_03996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04021_));
 sky130_fd_sc_hd__clkbuf_1 _09826_ (.A(_04021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[13] ));
 sky130_fd_sc_hd__and3_1 _09827_ (.A(_03939_),
    .B(_03893_),
    .C(_03988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04022_));
 sky130_fd_sc_hd__and2_1 _09828_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[14] ),
    .B(_04022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04023_));
 sky130_fd_sc_hd__nor2_1 _09829_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[14] ),
    .B(_04022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04024_));
 sky130_fd_sc_hd__or2_1 _09830_ (.A(_04023_),
    .B(_04024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04025_));
 sky130_fd_sc_hd__o21ba_1 _09831_ (.A1(_04007_),
    .A2(_04016_),
    .B1_N(_04017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04026_));
 sky130_fd_sc_hd__a41o_1 _09832_ (.A1(_04000_),
    .A2(_04010_),
    .A3(_04011_),
    .A4(_04018_),
    .B1(_04026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04027_));
 sky130_fd_sc_hd__xnor2_1 _09833_ (.A(_04025_),
    .B(_04027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04028_));
 sky130_fd_sc_hd__mux2_1 _09834_ (.A0(_04022_),
    .A1(_04028_),
    .S(_03996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04029_));
 sky130_fd_sc_hd__clkbuf_1 _09835_ (.A(_04029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[14] ));
 sky130_fd_sc_hd__and4_1 _09836_ (.A(_03939_),
    .B(_03935_),
    .C(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ),
    .D(_03988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04030_));
 sky130_fd_sc_hd__and2_1 _09837_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[15] ),
    .B(_04030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04031_));
 sky130_fd_sc_hd__nor2_1 _09838_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[15] ),
    .B(_04030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04032_));
 sky130_fd_sc_hd__nor2_1 _09839_ (.A(_04031_),
    .B(_04032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04033_));
 sky130_fd_sc_hd__inv_2 _09840_ (.A(_04025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04034_));
 sky130_fd_sc_hd__a21oi_1 _09841_ (.A1(_04034_),
    .A2(_04027_),
    .B1(_04023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04035_));
 sky130_fd_sc_hd__xnor2_1 _09842_ (.A(_04033_),
    .B(_04035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04036_));
 sky130_fd_sc_hd__mux2_1 _09843_ (.A0(_04030_),
    .A1(_04036_),
    .S(_03932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04037_));
 sky130_fd_sc_hd__clkbuf_1 _09844_ (.A(_04037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[15] ));
 sky130_fd_sc_hd__o21ba_1 _09845_ (.A1(_04023_),
    .A2(_04031_),
    .B1_N(_04032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04038_));
 sky130_fd_sc_hd__a31o_1 _09846_ (.A1(_04034_),
    .A2(_04027_),
    .A3(_04033_),
    .B1(_04038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04039_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09847_ (.A(_04039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04040_));
 sky130_fd_sc_hd__a21oi_1 _09848_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[16] ),
    .A2(_04040_),
    .B1(_03880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04041_));
 sky130_fd_sc_hd__o21a_1 _09849_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[16] ),
    .A2(_04040_),
    .B1(_04041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[16] ));
 sky130_fd_sc_hd__and2_1 _09850_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[16] ),
    .B(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04042_));
 sky130_fd_sc_hd__and2_1 _09851_ (.A(_04040_),
    .B(_04042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04043_));
 sky130_fd_sc_hd__a21o_1 _09852_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[16] ),
    .A2(_04040_),
    .B1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04044_));
 sky130_fd_sc_hd__and3b_1 _09853_ (.A_N(_04043_),
    .B(_03984_),
    .C(_04044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04045_));
 sky130_fd_sc_hd__clkbuf_1 _09854_ (.A(_04045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[17] ));
 sky130_fd_sc_hd__buf_2 _09855_ (.A(_03932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04046_));
 sky130_fd_sc_hd__o21ai_1 _09856_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[18] ),
    .A2(_04043_),
    .B1(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04047_));
 sky130_fd_sc_hd__a21oi_1 _09857_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[18] ),
    .A2(_04043_),
    .B1(_04047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[18] ));
 sky130_fd_sc_hd__and4_1 _09858_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[18] ),
    .B(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[19] ),
    .C(_04039_),
    .D(_04042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04048_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09859_ (.A(_04048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04049_));
 sky130_fd_sc_hd__a31o_1 _09860_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[18] ),
    .A2(_04040_),
    .A3(_04042_),
    .B1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04050_));
 sky130_fd_sc_hd__and3b_1 _09861_ (.A_N(_04049_),
    .B(_03984_),
    .C(_04050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04051_));
 sky130_fd_sc_hd__clkbuf_1 _09862_ (.A(_04051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[19] ));
 sky130_fd_sc_hd__and2_1 _09863_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[20] ),
    .B(_04049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04052_));
 sky130_fd_sc_hd__o21ai_1 _09864_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[20] ),
    .A2(_04049_),
    .B1(_03976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04053_));
 sky130_fd_sc_hd__nor2_1 _09865_ (.A(_04052_),
    .B(_04053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[20] ));
 sky130_fd_sc_hd__and2_1 _09866_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[20] ),
    .B(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04054_));
 sky130_fd_sc_hd__and2_1 _09867_ (.A(_04049_),
    .B(_04054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04055_));
 sky130_fd_sc_hd__inv_2 _09868_ (.A(_04055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04056_));
 sky130_fd_sc_hd__o211a_1 _09869_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[21] ),
    .A2(_04052_),
    .B1(_04056_),
    .C1(_03976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[21] ));
 sky130_fd_sc_hd__and3_1 _09870_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[22] ),
    .B(_04049_),
    .C(_04054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04057_));
 sky130_fd_sc_hd__o21ai_1 _09871_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[22] ),
    .A2(_04055_),
    .B1(_03976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04058_));
 sky130_fd_sc_hd__nor2_1 _09872_ (.A(_04057_),
    .B(_04058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[22] ));
 sky130_fd_sc_hd__and4_2 _09873_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[22] ),
    .B(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[23] ),
    .C(_04048_),
    .D(_04054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04059_));
 sky130_fd_sc_hd__o21ai_1 _09874_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[23] ),
    .A2(_04057_),
    .B1(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04060_));
 sky130_fd_sc_hd__nor2_1 _09875_ (.A(_04059_),
    .B(_04060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[23] ));
 sky130_fd_sc_hd__and2_1 _09876_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[24] ),
    .B(_04059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04061_));
 sky130_fd_sc_hd__o21ai_1 _09877_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[24] ),
    .A2(_04059_),
    .B1(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04062_));
 sky130_fd_sc_hd__nor2_1 _09878_ (.A(_04061_),
    .B(_04062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[24] ));
 sky130_fd_sc_hd__o21ai_1 _09879_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[25] ),
    .A2(_04061_),
    .B1(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04063_));
 sky130_fd_sc_hd__a21oi_1 _09880_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[25] ),
    .A2(_04061_),
    .B1(_04063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[25] ));
 sky130_fd_sc_hd__and4_1 _09881_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[24] ),
    .B(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[25] ),
    .C(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[26] ),
    .D(_04059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04064_));
 sky130_fd_sc_hd__a31o_1 _09882_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[24] ),
    .A2(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[25] ),
    .A3(_04059_),
    .B1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04065_));
 sky130_fd_sc_hd__and3b_1 _09883_ (.A_N(_04064_),
    .B(_03878_),
    .C(_04065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04066_));
 sky130_fd_sc_hd__clkbuf_1 _09884_ (.A(_04066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[26] ));
 sky130_fd_sc_hd__and2_1 _09885_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[27] ),
    .B(_04064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04067_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09886_ (.A(_04067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04068_));
 sky130_fd_sc_hd__o21ai_1 _09887_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[27] ),
    .A2(_04064_),
    .B1(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04069_));
 sky130_fd_sc_hd__nor2_1 _09888_ (.A(_04068_),
    .B(_04069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[27] ));
 sky130_fd_sc_hd__o21ai_1 _09889_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[28] ),
    .A2(_04068_),
    .B1(_03984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04070_));
 sky130_fd_sc_hd__a21oi_1 _09890_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[28] ),
    .A2(_04068_),
    .B1(_04070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[28] ));
 sky130_fd_sc_hd__a31o_1 _09891_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[27] ),
    .A2(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[28] ),
    .A3(_04064_),
    .B1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04071_));
 sky130_fd_sc_hd__and2_1 _09892_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[28] ),
    .B(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04072_));
 sky130_fd_sc_hd__nand2_1 _09893_ (.A(_04068_),
    .B(_04072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04073_));
 sky130_fd_sc_hd__and3_1 _09894_ (.A(_03984_),
    .B(_04071_),
    .C(_04073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04074_));
 sky130_fd_sc_hd__clkbuf_1 _09895_ (.A(_04074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[29] ));
 sky130_fd_sc_hd__inv_2 _09896_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04075_));
 sky130_fd_sc_hd__a31o_1 _09897_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[30] ),
    .A2(_04068_),
    .A3(_04072_),
    .B1(_03880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04076_));
 sky130_fd_sc_hd__a21oi_1 _09898_ (.A1(_04075_),
    .A2(_04073_),
    .B1(_04076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[30] ));
 sky130_fd_sc_hd__a41o_1 _09899_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[30] ),
    .A2(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[31] ),
    .A3(_04067_),
    .A4(_04072_),
    .B1(_03880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04077_));
 sky130_fd_sc_hd__a31o_1 _09900_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[30] ),
    .A2(_04067_),
    .A3(_04072_),
    .B1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04078_));
 sky130_fd_sc_hd__and2b_1 _09901_ (.A_N(_04077_),
    .B(_04078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04079_));
 sky130_fd_sc_hd__clkbuf_1 _09902_ (.A(_04079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[31] ));
 sky130_fd_sc_hd__clkbuf_4 _09903_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._01_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04080_));
 sky130_fd_sc_hd__clkbuf_2 _09904_ (.A(_04080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04081_));
 sky130_fd_sc_hd__mux2_1 _09905_ (.A0(\sa_inst.sak._23_[0] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[0] ),
    .S(_04081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04082_));
 sky130_fd_sc_hd__clkbuf_1 _09906_ (.A(_04082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ));
 sky130_fd_sc_hd__mux2_1 _09907_ (.A0(\sa_inst.sak._23_[1] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[1] ),
    .S(_04081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04083_));
 sky130_fd_sc_hd__clkbuf_1 _09908_ (.A(_04083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ));
 sky130_fd_sc_hd__mux2_1 _09909_ (.A0(\sa_inst.sak._23_[2] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[2] ),
    .S(_04081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04084_));
 sky130_fd_sc_hd__clkbuf_1 _09910_ (.A(_04084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ));
 sky130_fd_sc_hd__mux2_1 _09911_ (.A0(\sa_inst.sak._23_[3] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[3] ),
    .S(_04081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04085_));
 sky130_fd_sc_hd__clkbuf_1 _09912_ (.A(_04085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ));
 sky130_fd_sc_hd__mux2_1 _09913_ (.A0(\sa_inst.sak._23_[4] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[4] ),
    .S(_04081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04086_));
 sky130_fd_sc_hd__clkbuf_1 _09914_ (.A(_04086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ));
 sky130_fd_sc_hd__clkbuf_2 _09915_ (.A(_04080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04087_));
 sky130_fd_sc_hd__mux2_1 _09916_ (.A0(\sa_inst.sak._23_[5] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[5] ),
    .S(_04087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04088_));
 sky130_fd_sc_hd__clkbuf_1 _09917_ (.A(_04088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ));
 sky130_fd_sc_hd__mux2_1 _09918_ (.A0(\sa_inst.sak._23_[6] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[6] ),
    .S(_04087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04089_));
 sky130_fd_sc_hd__clkbuf_1 _09919_ (.A(_04089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ));
 sky130_fd_sc_hd__mux2_1 _09920_ (.A0(\sa_inst.sak._23_[7] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[7] ),
    .S(_04087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04090_));
 sky130_fd_sc_hd__clkbuf_1 _09921_ (.A(_04090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ));
 sky130_fd_sc_hd__mux2_1 _09922_ (.A0(\sa_inst.sak._23_[8] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[8] ),
    .S(_04087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04091_));
 sky130_fd_sc_hd__clkbuf_1 _09923_ (.A(_04091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ));
 sky130_fd_sc_hd__mux2_1 _09924_ (.A0(\sa_inst.sak._23_[9] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[9] ),
    .S(_04087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04092_));
 sky130_fd_sc_hd__clkbuf_1 _09925_ (.A(_04092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ));
 sky130_fd_sc_hd__clkbuf_2 _09926_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._01_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04093_));
 sky130_fd_sc_hd__mux2_1 _09927_ (.A0(\sa_inst.sak._23_[10] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[10] ),
    .S(_04093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04094_));
 sky130_fd_sc_hd__clkbuf_1 _09928_ (.A(_04094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ));
 sky130_fd_sc_hd__mux2_1 _09929_ (.A0(\sa_inst.sak._23_[11] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[11] ),
    .S(_04093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04095_));
 sky130_fd_sc_hd__clkbuf_1 _09930_ (.A(_04095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ));
 sky130_fd_sc_hd__mux2_1 _09931_ (.A0(\sa_inst.sak._23_[12] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[12] ),
    .S(_04093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04096_));
 sky130_fd_sc_hd__clkbuf_1 _09932_ (.A(_04096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ));
 sky130_fd_sc_hd__mux2_1 _09933_ (.A0(\sa_inst.sak._23_[13] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[13] ),
    .S(_04093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04097_));
 sky130_fd_sc_hd__clkbuf_1 _09934_ (.A(_04097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ));
 sky130_fd_sc_hd__mux2_1 _09935_ (.A0(\sa_inst.sak._23_[14] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[14] ),
    .S(_04093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04098_));
 sky130_fd_sc_hd__clkbuf_1 _09936_ (.A(_04098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ));
 sky130_fd_sc_hd__clkbuf_2 _09937_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._01_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04099_));
 sky130_fd_sc_hd__mux2_1 _09938_ (.A0(\sa_inst.sak._23_[15] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[15] ),
    .S(_04099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04100_));
 sky130_fd_sc_hd__clkbuf_1 _09939_ (.A(_04100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ));
 sky130_fd_sc_hd__mux2_1 _09940_ (.A0(\sa_inst.sak._23_[16] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[16] ),
    .S(_04099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04101_));
 sky130_fd_sc_hd__clkbuf_1 _09941_ (.A(_04101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ));
 sky130_fd_sc_hd__mux2_1 _09942_ (.A0(\sa_inst.sak._23_[17] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[17] ),
    .S(_04099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04102_));
 sky130_fd_sc_hd__clkbuf_1 _09943_ (.A(_04102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ));
 sky130_fd_sc_hd__mux2_1 _09944_ (.A0(\sa_inst.sak._23_[18] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[18] ),
    .S(_04099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04103_));
 sky130_fd_sc_hd__clkbuf_1 _09945_ (.A(_04103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ));
 sky130_fd_sc_hd__mux2_1 _09946_ (.A0(\sa_inst.sak._23_[19] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[19] ),
    .S(_04099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04104_));
 sky130_fd_sc_hd__clkbuf_1 _09947_ (.A(_04104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ));
 sky130_fd_sc_hd__clkbuf_2 _09948_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._01_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04105_));
 sky130_fd_sc_hd__mux2_1 _09949_ (.A0(\sa_inst.sak._23_[20] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[20] ),
    .S(_04105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04106_));
 sky130_fd_sc_hd__clkbuf_1 _09950_ (.A(_04106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ));
 sky130_fd_sc_hd__mux2_1 _09951_ (.A0(\sa_inst.sak._23_[21] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[21] ),
    .S(_04105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04107_));
 sky130_fd_sc_hd__clkbuf_1 _09952_ (.A(_04107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ));
 sky130_fd_sc_hd__mux2_1 _09953_ (.A0(\sa_inst.sak._23_[22] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[22] ),
    .S(_04105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04108_));
 sky130_fd_sc_hd__clkbuf_1 _09954_ (.A(_04108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ));
 sky130_fd_sc_hd__mux2_1 _09955_ (.A0(\sa_inst.sak._23_[23] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[23] ),
    .S(_04105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04109_));
 sky130_fd_sc_hd__clkbuf_1 _09956_ (.A(_04109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ));
 sky130_fd_sc_hd__mux2_1 _09957_ (.A0(\sa_inst.sak._23_[24] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[24] ),
    .S(_04105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04110_));
 sky130_fd_sc_hd__clkbuf_1 _09958_ (.A(_04110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ));
 sky130_fd_sc_hd__clkbuf_2 _09959_ (.A(\sa_inst.sak.rows:3.cols:3.pe_ij._01_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04111_));
 sky130_fd_sc_hd__mux2_1 _09960_ (.A0(\sa_inst.sak._23_[25] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[25] ),
    .S(_04111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04112_));
 sky130_fd_sc_hd__clkbuf_1 _09961_ (.A(_04112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ));
 sky130_fd_sc_hd__mux2_1 _09962_ (.A0(\sa_inst.sak._23_[26] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[26] ),
    .S(_04111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04113_));
 sky130_fd_sc_hd__clkbuf_1 _09963_ (.A(_04113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ));
 sky130_fd_sc_hd__mux2_1 _09964_ (.A0(\sa_inst.sak._23_[27] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[27] ),
    .S(_04111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04114_));
 sky130_fd_sc_hd__clkbuf_1 _09965_ (.A(_04114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ));
 sky130_fd_sc_hd__mux2_1 _09966_ (.A0(\sa_inst.sak._23_[28] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[28] ),
    .S(_04111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04115_));
 sky130_fd_sc_hd__clkbuf_1 _09967_ (.A(_04115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ));
 sky130_fd_sc_hd__mux2_1 _09968_ (.A0(\sa_inst.sak._23_[29] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[29] ),
    .S(_04111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04116_));
 sky130_fd_sc_hd__clkbuf_1 _09969_ (.A(_04116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ));
 sky130_fd_sc_hd__mux2_1 _09970_ (.A0(\sa_inst.sak._23_[30] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[30] ),
    .S(_04080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04117_));
 sky130_fd_sc_hd__clkbuf_1 _09971_ (.A(_04117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ));
 sky130_fd_sc_hd__mux2_1 _09972_ (.A0(\sa_inst.sak._23_[31] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[31] ),
    .S(_04080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04118_));
 sky130_fd_sc_hd__clkbuf_1 _09973_ (.A(_04118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ));
 sky130_fd_sc_hd__mux2_2 _09974_ (.A0(\sa_inst.sak._23_[32] ),
    .A1(\sa_inst.sak.rows:3.cols:3.pe_ij._02_ ),
    .S(_04080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04119_));
 sky130_fd_sc_hd__clkbuf_1 _09975_ (.A(_04119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ));
 sky130_fd_sc_hd__clkbuf_2 _09976_ (.A(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._10_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04120_));
 sky130_fd_sc_hd__and2b_1 _09977_ (.A_N(_04120_),
    .B(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04121_));
 sky130_fd_sc_hd__and2b_1 _09978_ (.A_N(_04120_),
    .B(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04122_));
 sky130_fd_sc_hd__mux2_1 _09979_ (.A0(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[5] ),
    .A1(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[3] ),
    .S(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._10_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04123_));
 sky130_fd_sc_hd__xnor2_1 _09980_ (.A(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._00_ ),
    .B(_04123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04124_));
 sky130_fd_sc_hd__clkbuf_2 _09981_ (.A(_04124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04125_));
 sky130_fd_sc_hd__mux2_1 _09982_ (.A0(_04121_),
    .A1(_04122_),
    .S(_04125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04126_));
 sky130_fd_sc_hd__clkbuf_1 _09983_ (.A(_04126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:2.a2s3_j._12_[1] ));
 sky130_fd_sc_hd__mux2_1 _09984_ (.A0(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[2] ),
    .A1(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[0] ),
    .S(_04120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04127_));
 sky130_fd_sc_hd__mux2_1 _09985_ (.A0(_04127_),
    .A1(_04121_),
    .S(_04125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04128_));
 sky130_fd_sc_hd__clkbuf_1 _09986_ (.A(_04128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:2.a2s3_j._12_[2] ));
 sky130_fd_sc_hd__mux2_1 _09987_ (.A0(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[3] ),
    .A1(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[1] ),
    .S(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._10_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04129_));
 sky130_fd_sc_hd__mux2_1 _09988_ (.A0(_04129_),
    .A1(_04127_),
    .S(_04125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04130_));
 sky130_fd_sc_hd__clkbuf_1 _09989_ (.A(_04130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:2.a2s3_j._12_[3] ));
 sky130_fd_sc_hd__mux2_1 _09990_ (.A0(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[4] ),
    .A1(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[2] ),
    .S(_04120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04131_));
 sky130_fd_sc_hd__mux2_1 _09991_ (.A0(_04131_),
    .A1(_04129_),
    .S(_04124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04132_));
 sky130_fd_sc_hd__clkbuf_1 _09992_ (.A(_04132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:2.a2s3_j._12_[4] ));
 sky130_fd_sc_hd__clkbuf_2 _09993_ (.A(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._10_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04133_));
 sky130_fd_sc_hd__and2b_1 _09994_ (.A_N(_04133_),
    .B(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04134_));
 sky130_fd_sc_hd__and2b_1 _09995_ (.A_N(_04133_),
    .B(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04135_));
 sky130_fd_sc_hd__mux2_1 _09996_ (.A0(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[5] ),
    .A1(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[3] ),
    .S(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._10_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04136_));
 sky130_fd_sc_hd__xnor2_1 _09997_ (.A(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._00_ ),
    .B(_04136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04137_));
 sky130_fd_sc_hd__clkbuf_2 _09998_ (.A(_04137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04138_));
 sky130_fd_sc_hd__mux2_1 _09999_ (.A0(_04134_),
    .A1(_04135_),
    .S(_04138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04139_));
 sky130_fd_sc_hd__clkbuf_1 _10000_ (.A(_04139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:1.a2s3_j._12_[1] ));
 sky130_fd_sc_hd__mux2_1 _10001_ (.A0(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[2] ),
    .A1(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[0] ),
    .S(_04133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04140_));
 sky130_fd_sc_hd__mux2_1 _10002_ (.A0(_04140_),
    .A1(_04134_),
    .S(_04138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04141_));
 sky130_fd_sc_hd__clkbuf_1 _10003_ (.A(_04141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:1.a2s3_j._12_[2] ));
 sky130_fd_sc_hd__mux2_1 _10004_ (.A0(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[3] ),
    .A1(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[1] ),
    .S(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._10_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04142_));
 sky130_fd_sc_hd__mux2_1 _10005_ (.A0(_04142_),
    .A1(_04140_),
    .S(_04138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04143_));
 sky130_fd_sc_hd__clkbuf_1 _10006_ (.A(_04143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:1.a2s3_j._12_[3] ));
 sky130_fd_sc_hd__mux2_1 _10007_ (.A0(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[4] ),
    .A1(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[2] ),
    .S(_04133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04144_));
 sky130_fd_sc_hd__mux2_1 _10008_ (.A0(_04144_),
    .A1(_04142_),
    .S(_04137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04145_));
 sky130_fd_sc_hd__clkbuf_1 _10009_ (.A(_04145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:1.a2s3_j._12_[4] ));
 sky130_fd_sc_hd__clkbuf_4 _10010_ (.A(\sa_inst.cols_l2a:3.l2a_i._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04146_));
 sky130_fd_sc_hd__xor2_2 _10011_ (.A(_04146_),
    .B(\sa_inst.cols_l2a:3.l2a_i._05_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04147_));
 sky130_fd_sc_hd__clkbuf_2 _10012_ (.A(_04147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._35_[0] ));
 sky130_fd_sc_hd__xor2_2 _10013_ (.A(_04146_),
    .B(\sa_inst.cols_l2a:3.l2a_i._05_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04148_));
 sky130_fd_sc_hd__clkbuf_2 _10014_ (.A(_04148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._35_[1] ));
 sky130_fd_sc_hd__xnor2_2 _10015_ (.A(_04146_),
    .B(\sa_inst.cols_l2a:3.l2a_i._05_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04149_));
 sky130_fd_sc_hd__inv_2 _10016_ (.A(_04149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:3.l2a_i._35_[2] ));
 sky130_fd_sc_hd__xnor2_2 _10017_ (.A(_04146_),
    .B(\sa_inst.cols_l2a:3.l2a_i._05_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04150_));
 sky130_fd_sc_hd__inv_2 _10018_ (.A(_04150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:3.l2a_i._35_[3] ));
 sky130_fd_sc_hd__inv_2 _10019_ (.A(_00830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:3.l2a_i._31_[0] ));
 sky130_fd_sc_hd__inv_2 _10020_ (.A(_00828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:3.l2a_i._31_[1] ));
 sky130_fd_sc_hd__a221o_1 _10021_ (.A1(\sa_inst.cols_l2a:3.l2a_i._31_[1] ),
    .A2(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._15_ ),
    .B1(\sa_inst.cols_l2a:3.l2a_i._31_[0] ),
    .B2(_00822_),
    .C1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._13_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._30_ ));
 sky130_fd_sc_hd__mux2_1 _10022_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[19] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[11] ),
    .S(_00848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04151_));
 sky130_fd_sc_hd__clkbuf_2 _10023_ (.A(_00848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04152_));
 sky130_fd_sc_hd__mux2_1 _10024_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[23] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[15] ),
    .S(_04152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04153_));
 sky130_fd_sc_hd__clkbuf_2 _10025_ (.A(_00847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04154_));
 sky130_fd_sc_hd__mux2_1 _10026_ (.A0(_04151_),
    .A1(_04153_),
    .S(_04154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04155_));
 sky130_fd_sc_hd__clkbuf_1 _10027_ (.A(_04155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[2] ));
 sky130_fd_sc_hd__mux2_1 _10028_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[20] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[12] ),
    .S(_04152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04156_));
 sky130_fd_sc_hd__mux2_1 _10029_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[24] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[16] ),
    .S(_04152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04157_));
 sky130_fd_sc_hd__mux2_1 _10030_ (.A0(_04156_),
    .A1(_04157_),
    .S(_04154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04158_));
 sky130_fd_sc_hd__clkbuf_1 _10031_ (.A(_04158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[3] ));
 sky130_fd_sc_hd__mux2_1 _10032_ (.A0(_00850_),
    .A1(_00971_),
    .S(_04154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04159_));
 sky130_fd_sc_hd__clkbuf_1 _10033_ (.A(_04159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[4] ));
 sky130_fd_sc_hd__mux2_1 _10034_ (.A0(_00853_),
    .A1(_00974_),
    .S(_00847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04160_));
 sky130_fd_sc_hd__clkbuf_1 _10035_ (.A(_04160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[5] ));
 sky130_fd_sc_hd__o22a_1 _10036_ (.A1(_00839_),
    .A2(_00845_),
    .B1(_04154_),
    .B2(_04153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[6] ));
 sky130_fd_sc_hd__a22o_1 _10037_ (.A1(_00840_),
    .A2(_00973_),
    .B1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._56_ ),
    .B2(_04157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[7] ));
 sky130_fd_sc_hd__mux2_1 _10038_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[17] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[1] ),
    .S(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._31_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04161_));
 sky130_fd_sc_hd__clkbuf_1 _10039_ (.A(_04161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[16] ));
 sky130_fd_sc_hd__mux2_1 _10040_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[18] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[2] ),
    .S(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._31_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04162_));
 sky130_fd_sc_hd__clkbuf_1 _10041_ (.A(_04162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[17] ));
 sky130_fd_sc_hd__mux2_1 _10042_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[19] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[3] ),
    .S(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._31_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04163_));
 sky130_fd_sc_hd__clkbuf_1 _10043_ (.A(_04163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[18] ));
 sky130_fd_sc_hd__mux2_1 _10044_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[20] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[4] ),
    .S(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._31_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04164_));
 sky130_fd_sc_hd__clkbuf_1 _10045_ (.A(_04164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[19] ));
 sky130_fd_sc_hd__mux2_1 _10046_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[21] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[5] ),
    .S(_00698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04165_));
 sky130_fd_sc_hd__clkbuf_1 _10047_ (.A(_04165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[20] ));
 sky130_fd_sc_hd__mux2_1 _10048_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[22] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[6] ),
    .S(_00698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04166_));
 sky130_fd_sc_hd__clkbuf_1 _10049_ (.A(_04166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[21] ));
 sky130_fd_sc_hd__mux2_1 _10050_ (.A0(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[23] ),
    .A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[7] ),
    .S(_00698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04167_));
 sky130_fd_sc_hd__clkbuf_1 _10051_ (.A(_04167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[22] ));
 sky130_fd_sc_hd__xnor2_1 _10052_ (.A(_04146_),
    .B(\sa_inst.cols_l2a:3.l2a_i._33_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04168_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10053_ (.A(_04168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._37_ ));
 sky130_fd_sc_hd__and2_1 _10054_ (.A(\sa_inst.cols_l2a:3.l2a_i._35_[3] ),
    .B(_04168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04169_));
 sky130_fd_sc_hd__a21o_1 _10055_ (.A1(\sa_inst.cols_l2a:3.l2a_i._02_[0] ),
    .A2(_04150_),
    .B1(_04169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.rshift._04_[0] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10056_ (.A(_04150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04170_));
 sky130_fd_sc_hd__a21o_1 _10057_ (.A1(\sa_inst.cols_l2a:3.l2a_i._02_[4] ),
    .A2(_04170_),
    .B1(_04169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04171_));
 sky130_fd_sc_hd__mux2_1 _10058_ (.A0(\sa_inst.cols_l2a:3.l2a_i.rshift._04_[0] ),
    .A1(_04171_),
    .S(\sa_inst.cols_l2a:3.l2a_i._35_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04172_));
 sky130_fd_sc_hd__clkbuf_1 _10059_ (.A(_04172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.rshift._10_[0] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10060_ (.A(_04169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04173_));
 sky130_fd_sc_hd__a21o_1 _10061_ (.A1(\sa_inst.cols_l2a:3.l2a_i._02_[2] ),
    .A2(_04170_),
    .B1(_04173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.rshift._04_[2] ));
 sky130_fd_sc_hd__nor2_1 _10062_ (.A(\sa_inst.cols_l2a:3.l2a_i._35_[3] ),
    .B(_04168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04174_));
 sky130_fd_sc_hd__or2_1 _10063_ (.A(_04173_),
    .B(_04174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04175_));
 sky130_fd_sc_hd__mux2_1 _10064_ (.A0(\sa_inst.cols_l2a:3.l2a_i.rshift._04_[2] ),
    .A1(_04175_),
    .S(\sa_inst.cols_l2a:3.l2a_i._35_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04176_));
 sky130_fd_sc_hd__mux2_1 _10065_ (.A0(\sa_inst.cols_l2a:3.l2a_i.rshift._10_[0] ),
    .A1(_04176_),
    .S(_04148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04177_));
 sky130_fd_sc_hd__clkbuf_1 _10066_ (.A(_04177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.rshift._17_[0] ));
 sky130_fd_sc_hd__a21o_1 _10067_ (.A1(\sa_inst.cols_l2a:3.l2a_i._02_[1] ),
    .A2(_04170_),
    .B1(_04173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.rshift._04_[1] ));
 sky130_fd_sc_hd__a21o_1 _10068_ (.A1(\sa_inst.cols_l2a:3.l2a_i._02_[5] ),
    .A2(_04170_),
    .B1(_04173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04178_));
 sky130_fd_sc_hd__mux2_1 _10069_ (.A0(\sa_inst.cols_l2a:3.l2a_i.rshift._04_[1] ),
    .A1(_04178_),
    .S(\sa_inst.cols_l2a:3.l2a_i._35_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04179_));
 sky130_fd_sc_hd__clkbuf_1 _10070_ (.A(_04179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.rshift._10_[1] ));
 sky130_fd_sc_hd__a21o_1 _10071_ (.A1(\sa_inst.cols_l2a:3.l2a_i._02_[3] ),
    .A2(_04170_),
    .B1(_04173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.rshift._04_[3] ));
 sky130_fd_sc_hd__and2_1 _10072_ (.A(\sa_inst.cols_l2a:3.l2a_i._35_[2] ),
    .B(\sa_inst.cols_l2a:3.l2a_i._37_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04180_));
 sky130_fd_sc_hd__a21o_1 _10073_ (.A1(_04149_),
    .A2(\sa_inst.cols_l2a:3.l2a_i.rshift._04_[3] ),
    .B1(_04180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04181_));
 sky130_fd_sc_hd__mux2_1 _10074_ (.A0(\sa_inst.cols_l2a:3.l2a_i.rshift._10_[1] ),
    .A1(_04181_),
    .S(\sa_inst.cols_l2a:3.l2a_i._35_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04182_));
 sky130_fd_sc_hd__mux2_1 _10075_ (.A0(\sa_inst.cols_l2a:3.l2a_i.rshift._17_[0] ),
    .A1(_04182_),
    .S(\sa_inst.cols_l2a:3.l2a_i._35_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04183_));
 sky130_fd_sc_hd__clkbuf_1 _10076_ (.A(_04183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._40_[0] ));
 sky130_fd_sc_hd__a21o_1 _10077_ (.A1(_04149_),
    .A2(_04171_),
    .B1(_04180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04184_));
 sky130_fd_sc_hd__mux2_1 _10078_ (.A0(_04176_),
    .A1(_04184_),
    .S(\sa_inst.cols_l2a:3.l2a_i._35_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04185_));
 sky130_fd_sc_hd__mux2_1 _10079_ (.A0(_04182_),
    .A1(_04185_),
    .S(\sa_inst.cols_l2a:3.l2a_i._35_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04186_));
 sky130_fd_sc_hd__clkbuf_1 _10080_ (.A(_04186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._40_[1] ));
 sky130_fd_sc_hd__a21o_1 _10081_ (.A1(_04149_),
    .A2(_04178_),
    .B1(_04180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04187_));
 sky130_fd_sc_hd__mux2_1 _10082_ (.A0(_04181_),
    .A1(_04187_),
    .S(\sa_inst.cols_l2a:3.l2a_i._35_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04188_));
 sky130_fd_sc_hd__mux2_1 _10083_ (.A0(_04185_),
    .A1(_04188_),
    .S(\sa_inst.cols_l2a:3.l2a_i._35_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04189_));
 sky130_fd_sc_hd__clkbuf_1 _10084_ (.A(_04189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._40_[2] ));
 sky130_fd_sc_hd__a21o_1 _10085_ (.A1(_04149_),
    .A2(_04175_),
    .B1(_04180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04190_));
 sky130_fd_sc_hd__mux2_1 _10086_ (.A0(_04184_),
    .A1(_04190_),
    .S(\sa_inst.cols_l2a:3.l2a_i._35_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04191_));
 sky130_fd_sc_hd__mux2_1 _10087_ (.A0(_04188_),
    .A1(_04191_),
    .S(\sa_inst.cols_l2a:3.l2a_i._35_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04192_));
 sky130_fd_sc_hd__clkbuf_1 _10088_ (.A(_04192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._40_[3] ));
 sky130_fd_sc_hd__mux2_1 _10089_ (.A0(_04187_),
    .A1(\sa_inst.cols_l2a:3.l2a_i._37_ ),
    .S(_04148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04193_));
 sky130_fd_sc_hd__mux2_1 _10090_ (.A0(_04191_),
    .A1(_04193_),
    .S(_04147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04194_));
 sky130_fd_sc_hd__clkbuf_1 _10091_ (.A(_04194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._40_[4] ));
 sky130_fd_sc_hd__mux2_1 _10092_ (.A0(_04190_),
    .A1(\sa_inst.cols_l2a:3.l2a_i._37_ ),
    .S(_04148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04195_));
 sky130_fd_sc_hd__mux2_1 _10093_ (.A0(_04193_),
    .A1(_04195_),
    .S(_04147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04196_));
 sky130_fd_sc_hd__clkbuf_1 _10094_ (.A(_04196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._40_[5] ));
 sky130_fd_sc_hd__mux2_1 _10095_ (.A0(_04195_),
    .A1(\sa_inst.cols_l2a:3.l2a_i._37_ ),
    .S(_04147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04197_));
 sky130_fd_sc_hd__clkbuf_1 _10096_ (.A(_04197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._40_[6] ));
 sky130_fd_sc_hd__clkbuf_4 _10097_ (.A(\sa_inst.cols_l2a:2.l2a_i._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04198_));
 sky130_fd_sc_hd__xor2_2 _10098_ (.A(_04198_),
    .B(\sa_inst.cols_l2a:2.l2a_i._05_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04199_));
 sky130_fd_sc_hd__clkbuf_2 _10099_ (.A(_04199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._35_[0] ));
 sky130_fd_sc_hd__xor2_2 _10100_ (.A(_04198_),
    .B(\sa_inst.cols_l2a:2.l2a_i._05_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04200_));
 sky130_fd_sc_hd__clkbuf_2 _10101_ (.A(_04200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._35_[1] ));
 sky130_fd_sc_hd__xnor2_2 _10102_ (.A(_04198_),
    .B(\sa_inst.cols_l2a:2.l2a_i._05_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04201_));
 sky130_fd_sc_hd__inv_2 _10103_ (.A(_04201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:2.l2a_i._35_[2] ));
 sky130_fd_sc_hd__xnor2_1 _10104_ (.A(_04198_),
    .B(\sa_inst.cols_l2a:2.l2a_i._05_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04202_));
 sky130_fd_sc_hd__inv_2 _10105_ (.A(_04202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:2.l2a_i._35_[3] ));
 sky130_fd_sc_hd__inv_2 _10106_ (.A(_00880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:2.l2a_i._31_[0] ));
 sky130_fd_sc_hd__inv_2 _10107_ (.A(_00878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:2.l2a_i._31_[1] ));
 sky130_fd_sc_hd__a221o_1 _10108_ (.A1(\sa_inst.cols_l2a:2.l2a_i._31_[1] ),
    .A2(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._15_ ),
    .B1(\sa_inst.cols_l2a:2.l2a_i._31_[0] ),
    .B2(_00872_),
    .C1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._13_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._30_ ));
 sky130_fd_sc_hd__mux2_1 _10109_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[19] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[11] ),
    .S(_00898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04203_));
 sky130_fd_sc_hd__clkbuf_2 _10110_ (.A(_00898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04204_));
 sky130_fd_sc_hd__mux2_1 _10111_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[23] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[15] ),
    .S(_04204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04205_));
 sky130_fd_sc_hd__clkbuf_2 _10112_ (.A(_00897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04206_));
 sky130_fd_sc_hd__mux2_1 _10113_ (.A0(_04203_),
    .A1(_04205_),
    .S(_04206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04207_));
 sky130_fd_sc_hd__clkbuf_1 _10114_ (.A(_04207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[2] ));
 sky130_fd_sc_hd__mux2_1 _10115_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[20] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[12] ),
    .S(_04204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04208_));
 sky130_fd_sc_hd__mux2_1 _10116_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[24] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[16] ),
    .S(_04204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04209_));
 sky130_fd_sc_hd__mux2_1 _10117_ (.A0(_04208_),
    .A1(_04209_),
    .S(_04206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04210_));
 sky130_fd_sc_hd__clkbuf_1 _10118_ (.A(_04210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[3] ));
 sky130_fd_sc_hd__mux2_1 _10119_ (.A0(_00900_),
    .A1(_00992_),
    .S(_04206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04211_));
 sky130_fd_sc_hd__clkbuf_1 _10120_ (.A(_04211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[4] ));
 sky130_fd_sc_hd__mux2_1 _10121_ (.A0(_00903_),
    .A1(_00995_),
    .S(_00897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04212_));
 sky130_fd_sc_hd__clkbuf_1 _10122_ (.A(_04212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[5] ));
 sky130_fd_sc_hd__o22a_1 _10123_ (.A1(_00889_),
    .A2(_00895_),
    .B1(_04206_),
    .B2(_04205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[6] ));
 sky130_fd_sc_hd__a22o_1 _10124_ (.A1(_00890_),
    .A2(_00994_),
    .B1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._56_ ),
    .B2(_04209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[7] ));
 sky130_fd_sc_hd__mux2_1 _10125_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[17] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[1] ),
    .S(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._31_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04213_));
 sky130_fd_sc_hd__clkbuf_1 _10126_ (.A(_04213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[16] ));
 sky130_fd_sc_hd__mux2_1 _10127_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[18] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[2] ),
    .S(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._31_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04214_));
 sky130_fd_sc_hd__clkbuf_1 _10128_ (.A(_04214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[17] ));
 sky130_fd_sc_hd__mux2_1 _10129_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[19] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[3] ),
    .S(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._31_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04215_));
 sky130_fd_sc_hd__clkbuf_1 _10130_ (.A(_04215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[18] ));
 sky130_fd_sc_hd__mux2_1 _10131_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[20] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[4] ),
    .S(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._31_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04216_));
 sky130_fd_sc_hd__clkbuf_1 _10132_ (.A(_04216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[19] ));
 sky130_fd_sc_hd__mux2_1 _10133_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[21] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[5] ),
    .S(_00738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04217_));
 sky130_fd_sc_hd__clkbuf_1 _10134_ (.A(_04217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[20] ));
 sky130_fd_sc_hd__mux2_1 _10135_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[22] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[6] ),
    .S(_00738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04218_));
 sky130_fd_sc_hd__clkbuf_1 _10136_ (.A(_04218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[21] ));
 sky130_fd_sc_hd__mux2_1 _10137_ (.A0(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[23] ),
    .A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[7] ),
    .S(_00738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04219_));
 sky130_fd_sc_hd__clkbuf_1 _10138_ (.A(_04219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[22] ));
 sky130_fd_sc_hd__xnor2_1 _10139_ (.A(_04198_),
    .B(\sa_inst.cols_l2a:2.l2a_i._33_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04220_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10140_ (.A(_04220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._37_ ));
 sky130_fd_sc_hd__and2_1 _10141_ (.A(\sa_inst.cols_l2a:2.l2a_i._35_[3] ),
    .B(_04220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04221_));
 sky130_fd_sc_hd__a21o_1 _10142_ (.A1(\sa_inst.cols_l2a:2.l2a_i._02_[0] ),
    .A2(_04202_),
    .B1(_04221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.rshift._04_[0] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10143_ (.A(_04202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04222_));
 sky130_fd_sc_hd__a21o_1 _10144_ (.A1(\sa_inst.cols_l2a:2.l2a_i._02_[4] ),
    .A2(_04222_),
    .B1(_04221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04223_));
 sky130_fd_sc_hd__mux2_1 _10145_ (.A0(\sa_inst.cols_l2a:2.l2a_i.rshift._04_[0] ),
    .A1(_04223_),
    .S(\sa_inst.cols_l2a:2.l2a_i._35_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04224_));
 sky130_fd_sc_hd__clkbuf_1 _10146_ (.A(_04224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.rshift._10_[0] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10147_ (.A(_04221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04225_));
 sky130_fd_sc_hd__a21o_1 _10148_ (.A1(\sa_inst.cols_l2a:2.l2a_i._02_[2] ),
    .A2(_04222_),
    .B1(_04225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.rshift._04_[2] ));
 sky130_fd_sc_hd__nor2_1 _10149_ (.A(\sa_inst.cols_l2a:2.l2a_i._35_[3] ),
    .B(_04220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04226_));
 sky130_fd_sc_hd__or2_1 _10150_ (.A(_04225_),
    .B(_04226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04227_));
 sky130_fd_sc_hd__mux2_1 _10151_ (.A0(\sa_inst.cols_l2a:2.l2a_i.rshift._04_[2] ),
    .A1(_04227_),
    .S(\sa_inst.cols_l2a:2.l2a_i._35_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04228_));
 sky130_fd_sc_hd__mux2_1 _10152_ (.A0(\sa_inst.cols_l2a:2.l2a_i.rshift._10_[0] ),
    .A1(_04228_),
    .S(_04200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04229_));
 sky130_fd_sc_hd__clkbuf_1 _10153_ (.A(_04229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.rshift._17_[0] ));
 sky130_fd_sc_hd__a21o_1 _10154_ (.A1(\sa_inst.cols_l2a:2.l2a_i._02_[1] ),
    .A2(_04222_),
    .B1(_04225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.rshift._04_[1] ));
 sky130_fd_sc_hd__a21o_1 _10155_ (.A1(\sa_inst.cols_l2a:2.l2a_i._02_[5] ),
    .A2(_04222_),
    .B1(_04225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04230_));
 sky130_fd_sc_hd__mux2_1 _10156_ (.A0(\sa_inst.cols_l2a:2.l2a_i.rshift._04_[1] ),
    .A1(_04230_),
    .S(\sa_inst.cols_l2a:2.l2a_i._35_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04231_));
 sky130_fd_sc_hd__clkbuf_1 _10157_ (.A(_04231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.rshift._10_[1] ));
 sky130_fd_sc_hd__a21o_1 _10158_ (.A1(\sa_inst.cols_l2a:2.l2a_i._02_[3] ),
    .A2(_04222_),
    .B1(_04225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.rshift._04_[3] ));
 sky130_fd_sc_hd__and2_1 _10159_ (.A(\sa_inst.cols_l2a:2.l2a_i._35_[2] ),
    .B(\sa_inst.cols_l2a:2.l2a_i._37_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04232_));
 sky130_fd_sc_hd__a21o_1 _10160_ (.A1(_04201_),
    .A2(\sa_inst.cols_l2a:2.l2a_i.rshift._04_[3] ),
    .B1(_04232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04233_));
 sky130_fd_sc_hd__mux2_1 _10161_ (.A0(\sa_inst.cols_l2a:2.l2a_i.rshift._10_[1] ),
    .A1(_04233_),
    .S(\sa_inst.cols_l2a:2.l2a_i._35_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04234_));
 sky130_fd_sc_hd__mux2_1 _10162_ (.A0(\sa_inst.cols_l2a:2.l2a_i.rshift._17_[0] ),
    .A1(_04234_),
    .S(\sa_inst.cols_l2a:2.l2a_i._35_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04235_));
 sky130_fd_sc_hd__clkbuf_1 _10163_ (.A(_04235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._40_[0] ));
 sky130_fd_sc_hd__a21o_1 _10164_ (.A1(_04201_),
    .A2(_04223_),
    .B1(_04232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04236_));
 sky130_fd_sc_hd__mux2_1 _10165_ (.A0(_04228_),
    .A1(_04236_),
    .S(\sa_inst.cols_l2a:2.l2a_i._35_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04237_));
 sky130_fd_sc_hd__mux2_1 _10166_ (.A0(_04234_),
    .A1(_04237_),
    .S(\sa_inst.cols_l2a:2.l2a_i._35_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04238_));
 sky130_fd_sc_hd__clkbuf_1 _10167_ (.A(_04238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._40_[1] ));
 sky130_fd_sc_hd__a21o_1 _10168_ (.A1(_04201_),
    .A2(_04230_),
    .B1(_04232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04239_));
 sky130_fd_sc_hd__mux2_1 _10169_ (.A0(_04233_),
    .A1(_04239_),
    .S(\sa_inst.cols_l2a:2.l2a_i._35_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04240_));
 sky130_fd_sc_hd__mux2_1 _10170_ (.A0(_04237_),
    .A1(_04240_),
    .S(\sa_inst.cols_l2a:2.l2a_i._35_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04241_));
 sky130_fd_sc_hd__clkbuf_1 _10171_ (.A(_04241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._40_[2] ));
 sky130_fd_sc_hd__a21o_1 _10172_ (.A1(_04201_),
    .A2(_04227_),
    .B1(_04232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04242_));
 sky130_fd_sc_hd__mux2_1 _10173_ (.A0(_04236_),
    .A1(_04242_),
    .S(\sa_inst.cols_l2a:2.l2a_i._35_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04243_));
 sky130_fd_sc_hd__mux2_1 _10174_ (.A0(_04240_),
    .A1(_04243_),
    .S(\sa_inst.cols_l2a:2.l2a_i._35_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04244_));
 sky130_fd_sc_hd__clkbuf_1 _10175_ (.A(_04244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._40_[3] ));
 sky130_fd_sc_hd__mux2_1 _10176_ (.A0(_04239_),
    .A1(\sa_inst.cols_l2a:2.l2a_i._37_ ),
    .S(_04200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04245_));
 sky130_fd_sc_hd__mux2_1 _10177_ (.A0(_04243_),
    .A1(_04245_),
    .S(_04199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04246_));
 sky130_fd_sc_hd__clkbuf_1 _10178_ (.A(_04246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._40_[4] ));
 sky130_fd_sc_hd__mux2_1 _10179_ (.A0(_04242_),
    .A1(\sa_inst.cols_l2a:2.l2a_i._37_ ),
    .S(_04200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04247_));
 sky130_fd_sc_hd__mux2_1 _10180_ (.A0(_04245_),
    .A1(_04247_),
    .S(_04199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04248_));
 sky130_fd_sc_hd__clkbuf_1 _10181_ (.A(_04248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._40_[5] ));
 sky130_fd_sc_hd__mux2_1 _10182_ (.A0(_04247_),
    .A1(\sa_inst.cols_l2a:2.l2a_i._37_ ),
    .S(_04199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04249_));
 sky130_fd_sc_hd__clkbuf_1 _10183_ (.A(_04249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._40_[6] ));
 sky130_fd_sc_hd__clkbuf_4 _10184_ (.A(\sa_inst.cols_l2a:1.l2a_i._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04250_));
 sky130_fd_sc_hd__xor2_2 _10185_ (.A(_04250_),
    .B(\sa_inst.cols_l2a:1.l2a_i._05_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04251_));
 sky130_fd_sc_hd__clkbuf_2 _10186_ (.A(_04251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._35_[0] ));
 sky130_fd_sc_hd__xor2_2 _10187_ (.A(_04250_),
    .B(\sa_inst.cols_l2a:1.l2a_i._05_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04252_));
 sky130_fd_sc_hd__clkbuf_2 _10188_ (.A(_04252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._35_[1] ));
 sky130_fd_sc_hd__xnor2_2 _10189_ (.A(_04250_),
    .B(\sa_inst.cols_l2a:1.l2a_i._05_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04253_));
 sky130_fd_sc_hd__inv_2 _10190_ (.A(_04253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:1.l2a_i._35_[2] ));
 sky130_fd_sc_hd__xnor2_1 _10191_ (.A(_04250_),
    .B(\sa_inst.cols_l2a:1.l2a_i._05_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04254_));
 sky130_fd_sc_hd__inv_2 _10192_ (.A(_04254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:1.l2a_i._35_[3] ));
 sky130_fd_sc_hd__inv_2 _10193_ (.A(_00930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:1.l2a_i._31_[0] ));
 sky130_fd_sc_hd__inv_2 _10194_ (.A(_00928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:1.l2a_i._31_[1] ));
 sky130_fd_sc_hd__a221o_1 _10195_ (.A1(\sa_inst.cols_l2a:1.l2a_i._31_[1] ),
    .A2(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._15_ ),
    .B1(\sa_inst.cols_l2a:1.l2a_i._31_[0] ),
    .B2(_00922_),
    .C1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._13_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._30_ ));
 sky130_fd_sc_hd__mux2_1 _10196_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[19] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[11] ),
    .S(_00948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04255_));
 sky130_fd_sc_hd__clkbuf_2 _10197_ (.A(_00948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04256_));
 sky130_fd_sc_hd__mux2_1 _10198_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[23] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[15] ),
    .S(_04256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04257_));
 sky130_fd_sc_hd__clkbuf_2 _10199_ (.A(_00947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04258_));
 sky130_fd_sc_hd__mux2_1 _10200_ (.A0(_04255_),
    .A1(_04257_),
    .S(_04258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04259_));
 sky130_fd_sc_hd__clkbuf_1 _10201_ (.A(_04259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[2] ));
 sky130_fd_sc_hd__mux2_1 _10202_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[20] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[12] ),
    .S(_04256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04260_));
 sky130_fd_sc_hd__mux2_1 _10203_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[24] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[16] ),
    .S(_04256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04261_));
 sky130_fd_sc_hd__mux2_1 _10204_ (.A0(_04260_),
    .A1(_04261_),
    .S(_04258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04262_));
 sky130_fd_sc_hd__clkbuf_1 _10205_ (.A(_04262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[3] ));
 sky130_fd_sc_hd__mux2_1 _10206_ (.A0(_00950_),
    .A1(_01012_),
    .S(_04258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04263_));
 sky130_fd_sc_hd__clkbuf_1 _10207_ (.A(_04263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[4] ));
 sky130_fd_sc_hd__mux2_1 _10208_ (.A0(_00953_),
    .A1(_01015_),
    .S(_00947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04264_));
 sky130_fd_sc_hd__clkbuf_1 _10209_ (.A(_04264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[5] ));
 sky130_fd_sc_hd__o22a_1 _10210_ (.A1(_00939_),
    .A2(_00945_),
    .B1(_04258_),
    .B2(_04257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[6] ));
 sky130_fd_sc_hd__a22o_1 _10211_ (.A1(_00940_),
    .A2(_01014_),
    .B1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._56_ ),
    .B2(_04261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[7] ));
 sky130_fd_sc_hd__mux2_1 _10212_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[17] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[1] ),
    .S(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._31_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04265_));
 sky130_fd_sc_hd__clkbuf_1 _10213_ (.A(_04265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[16] ));
 sky130_fd_sc_hd__mux2_1 _10214_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[18] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[2] ),
    .S(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._31_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04266_));
 sky130_fd_sc_hd__clkbuf_1 _10215_ (.A(_04266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[17] ));
 sky130_fd_sc_hd__mux2_1 _10216_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[19] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[3] ),
    .S(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._31_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04267_));
 sky130_fd_sc_hd__clkbuf_1 _10217_ (.A(_04267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[18] ));
 sky130_fd_sc_hd__mux2_1 _10218_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[20] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[4] ),
    .S(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._31_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04268_));
 sky130_fd_sc_hd__clkbuf_1 _10219_ (.A(_04268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[19] ));
 sky130_fd_sc_hd__mux2_1 _10220_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[21] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[5] ),
    .S(_00778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04269_));
 sky130_fd_sc_hd__clkbuf_1 _10221_ (.A(_04269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[20] ));
 sky130_fd_sc_hd__mux2_1 _10222_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[22] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[6] ),
    .S(_00778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04270_));
 sky130_fd_sc_hd__clkbuf_1 _10223_ (.A(_04270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[21] ));
 sky130_fd_sc_hd__mux2_1 _10224_ (.A0(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[23] ),
    .A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[7] ),
    .S(_00778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04271_));
 sky130_fd_sc_hd__clkbuf_1 _10225_ (.A(_04271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[22] ));
 sky130_fd_sc_hd__xnor2_1 _10226_ (.A(_04250_),
    .B(\sa_inst.cols_l2a:1.l2a_i._33_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04272_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10227_ (.A(_04272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._37_ ));
 sky130_fd_sc_hd__and2_1 _10228_ (.A(\sa_inst.cols_l2a:1.l2a_i._35_[3] ),
    .B(_04272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04273_));
 sky130_fd_sc_hd__a21o_1 _10229_ (.A1(\sa_inst.cols_l2a:1.l2a_i._02_[0] ),
    .A2(_04254_),
    .B1(_04273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.rshift._04_[0] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10230_ (.A(_04254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04274_));
 sky130_fd_sc_hd__a21o_1 _10231_ (.A1(\sa_inst.cols_l2a:1.l2a_i._02_[4] ),
    .A2(_04274_),
    .B1(_04273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04275_));
 sky130_fd_sc_hd__mux2_1 _10232_ (.A0(\sa_inst.cols_l2a:1.l2a_i.rshift._04_[0] ),
    .A1(_04275_),
    .S(\sa_inst.cols_l2a:1.l2a_i._35_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04276_));
 sky130_fd_sc_hd__clkbuf_1 _10233_ (.A(_04276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.rshift._10_[0] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10234_ (.A(_04273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04277_));
 sky130_fd_sc_hd__a21o_1 _10235_ (.A1(\sa_inst.cols_l2a:1.l2a_i._02_[2] ),
    .A2(_04274_),
    .B1(_04277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.rshift._04_[2] ));
 sky130_fd_sc_hd__nor2_1 _10236_ (.A(\sa_inst.cols_l2a:1.l2a_i._35_[3] ),
    .B(_04272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04278_));
 sky130_fd_sc_hd__or2_1 _10237_ (.A(_04277_),
    .B(_04278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04279_));
 sky130_fd_sc_hd__mux2_1 _10238_ (.A0(\sa_inst.cols_l2a:1.l2a_i.rshift._04_[2] ),
    .A1(_04279_),
    .S(\sa_inst.cols_l2a:1.l2a_i._35_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04280_));
 sky130_fd_sc_hd__mux2_1 _10239_ (.A0(\sa_inst.cols_l2a:1.l2a_i.rshift._10_[0] ),
    .A1(_04280_),
    .S(_04252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04281_));
 sky130_fd_sc_hd__clkbuf_1 _10240_ (.A(_04281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.rshift._17_[0] ));
 sky130_fd_sc_hd__a21o_1 _10241_ (.A1(\sa_inst.cols_l2a:1.l2a_i._02_[1] ),
    .A2(_04274_),
    .B1(_04277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.rshift._04_[1] ));
 sky130_fd_sc_hd__a21o_1 _10242_ (.A1(\sa_inst.cols_l2a:1.l2a_i._02_[5] ),
    .A2(_04274_),
    .B1(_04277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04282_));
 sky130_fd_sc_hd__mux2_1 _10243_ (.A0(\sa_inst.cols_l2a:1.l2a_i.rshift._04_[1] ),
    .A1(_04282_),
    .S(\sa_inst.cols_l2a:1.l2a_i._35_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04283_));
 sky130_fd_sc_hd__clkbuf_1 _10244_ (.A(_04283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.rshift._10_[1] ));
 sky130_fd_sc_hd__a21o_1 _10245_ (.A1(\sa_inst.cols_l2a:1.l2a_i._02_[3] ),
    .A2(_04274_),
    .B1(_04277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.rshift._04_[3] ));
 sky130_fd_sc_hd__and2_1 _10246_ (.A(\sa_inst.cols_l2a:1.l2a_i._35_[2] ),
    .B(\sa_inst.cols_l2a:1.l2a_i._37_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04284_));
 sky130_fd_sc_hd__a21o_1 _10247_ (.A1(_04253_),
    .A2(\sa_inst.cols_l2a:1.l2a_i.rshift._04_[3] ),
    .B1(_04284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04285_));
 sky130_fd_sc_hd__mux2_1 _10248_ (.A0(\sa_inst.cols_l2a:1.l2a_i.rshift._10_[1] ),
    .A1(_04285_),
    .S(\sa_inst.cols_l2a:1.l2a_i._35_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04286_));
 sky130_fd_sc_hd__mux2_1 _10249_ (.A0(\sa_inst.cols_l2a:1.l2a_i.rshift._17_[0] ),
    .A1(_04286_),
    .S(\sa_inst.cols_l2a:1.l2a_i._35_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04287_));
 sky130_fd_sc_hd__clkbuf_1 _10250_ (.A(_04287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._40_[0] ));
 sky130_fd_sc_hd__a21o_1 _10251_ (.A1(_04253_),
    .A2(_04275_),
    .B1(_04284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04288_));
 sky130_fd_sc_hd__mux2_1 _10252_ (.A0(_04280_),
    .A1(_04288_),
    .S(\sa_inst.cols_l2a:1.l2a_i._35_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04289_));
 sky130_fd_sc_hd__mux2_1 _10253_ (.A0(_04286_),
    .A1(_04289_),
    .S(\sa_inst.cols_l2a:1.l2a_i._35_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04290_));
 sky130_fd_sc_hd__clkbuf_1 _10254_ (.A(_04290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._40_[1] ));
 sky130_fd_sc_hd__a21o_1 _10255_ (.A1(_04253_),
    .A2(_04282_),
    .B1(_04284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04291_));
 sky130_fd_sc_hd__mux2_1 _10256_ (.A0(_04285_),
    .A1(_04291_),
    .S(\sa_inst.cols_l2a:1.l2a_i._35_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04292_));
 sky130_fd_sc_hd__mux2_1 _10257_ (.A0(_04289_),
    .A1(_04292_),
    .S(\sa_inst.cols_l2a:1.l2a_i._35_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04293_));
 sky130_fd_sc_hd__clkbuf_1 _10258_ (.A(_04293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._40_[2] ));
 sky130_fd_sc_hd__a21o_1 _10259_ (.A1(_04253_),
    .A2(_04279_),
    .B1(_04284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04294_));
 sky130_fd_sc_hd__mux2_1 _10260_ (.A0(_04288_),
    .A1(_04294_),
    .S(\sa_inst.cols_l2a:1.l2a_i._35_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04295_));
 sky130_fd_sc_hd__mux2_1 _10261_ (.A0(_04292_),
    .A1(_04295_),
    .S(\sa_inst.cols_l2a:1.l2a_i._35_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04296_));
 sky130_fd_sc_hd__clkbuf_1 _10262_ (.A(_04296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._40_[3] ));
 sky130_fd_sc_hd__mux2_1 _10263_ (.A0(_04291_),
    .A1(\sa_inst.cols_l2a:1.l2a_i._37_ ),
    .S(_04252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04297_));
 sky130_fd_sc_hd__mux2_1 _10264_ (.A0(_04295_),
    .A1(_04297_),
    .S(_04251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04298_));
 sky130_fd_sc_hd__clkbuf_1 _10265_ (.A(_04298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._40_[4] ));
 sky130_fd_sc_hd__mux2_1 _10266_ (.A0(_04294_),
    .A1(\sa_inst.cols_l2a:1.l2a_i._37_ ),
    .S(_04252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04299_));
 sky130_fd_sc_hd__mux2_1 _10267_ (.A0(_04297_),
    .A1(_04299_),
    .S(_04251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04300_));
 sky130_fd_sc_hd__clkbuf_1 _10268_ (.A(_04300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._40_[5] ));
 sky130_fd_sc_hd__mux2_1 _10269_ (.A0(_04299_),
    .A1(\sa_inst.cols_l2a:1.l2a_i._37_ ),
    .S(_04251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04301_));
 sky130_fd_sc_hd__clkbuf_1 _10270_ (.A(_04301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._40_[6] ));
 sky130_fd_sc_hd__clkbuf_2 _10271_ (.A(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._10_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04302_));
 sky130_fd_sc_hd__and2b_1 _10272_ (.A_N(_04302_),
    .B(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04303_));
 sky130_fd_sc_hd__and2b_1 _10273_ (.A_N(_04302_),
    .B(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04304_));
 sky130_fd_sc_hd__mux2_1 _10274_ (.A0(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[5] ),
    .A1(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[3] ),
    .S(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._10_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04305_));
 sky130_fd_sc_hd__xnor2_1 _10275_ (.A(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._00_ ),
    .B(_04305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04306_));
 sky130_fd_sc_hd__clkbuf_2 _10276_ (.A(_04306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04307_));
 sky130_fd_sc_hd__mux2_1 _10277_ (.A0(_04303_),
    .A1(_04304_),
    .S(_04307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04308_));
 sky130_fd_sc_hd__clkbuf_1 _10278_ (.A(_04308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:3.a2s3_j._12_[1] ));
 sky130_fd_sc_hd__mux2_1 _10279_ (.A0(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[2] ),
    .A1(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[0] ),
    .S(_04302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04309_));
 sky130_fd_sc_hd__mux2_1 _10280_ (.A0(_04309_),
    .A1(_04303_),
    .S(_04307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04310_));
 sky130_fd_sc_hd__clkbuf_1 _10281_ (.A(_04310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:3.a2s3_j._12_[2] ));
 sky130_fd_sc_hd__mux2_1 _10282_ (.A0(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[3] ),
    .A1(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[1] ),
    .S(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._10_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04311_));
 sky130_fd_sc_hd__mux2_1 _10283_ (.A0(_04311_),
    .A1(_04309_),
    .S(_04307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04312_));
 sky130_fd_sc_hd__clkbuf_1 _10284_ (.A(_04312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:3.a2s3_j._12_[3] ));
 sky130_fd_sc_hd__mux2_1 _10285_ (.A0(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[4] ),
    .A1(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[2] ),
    .S(_04302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04313_));
 sky130_fd_sc_hd__mux2_1 _10286_ (.A0(_04313_),
    .A1(_04311_),
    .S(_04306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04314_));
 sky130_fd_sc_hd__clkbuf_1 _10287_ (.A(_04314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:3.a2s3_j._12_[4] ));
 sky130_fd_sc_hd__inv_2 _10288_ (.A(\sa_inst._22_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._17_ ));
 sky130_fd_sc_hd__clkinv_2 _10289_ (.A(\sa_inst.sak._22_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._17_ ));
 sky130_fd_sc_hd__clkinv_2 _10290_ (.A(\sa_inst.sak._09_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._17_ ));
 sky130_fd_sc_hd__clkinv_2 _10291_ (.A(\sa_inst.sak._04_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._17_ ));
 sky130_fd_sc_hd__clkinv_2 _10292_ (.A(\sa_inst.sak._20_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._17_ ));
 sky130_fd_sc_hd__clkbuf_1 _10293_ (.A(_00813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04315_));
 sky130_fd_sc_hd__o21ai_1 _10294_ (.A1(net1),
    .A2(net12),
    .B1(_04315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04316_));
 sky130_fd_sc_hd__nand3_1 _10295_ (.A(_00817_),
    .B(_01045_),
    .C(_04316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_a2s3:1.a2s3_j._07_ ));
 sky130_fd_sc_hd__or2_1 _10296_ (.A(net23),
    .B(_01045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04317_));
 sky130_fd_sc_hd__o21a_1 _10297_ (.A1(net24),
    .A2(_00814_),
    .B1(_04317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:1.a2s3_j._14_[0] ));
 sky130_fd_sc_hd__or4_1 _10298_ (.A(\sa_inst._17_[0] ),
    .B(\sa_inst._17_[1] ),
    .C(\sa_inst._17_[7] ),
    .D(_00806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04318_));
 sky130_fd_sc_hd__clkbuf_1 _10299_ (.A(_04318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:3.a2s3_j._07_ ));
 sky130_fd_sc_hd__xnor2_1 _10300_ (.A(\sa_inst._17_[6] ),
    .B(\sa_inst._17_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_a2s3:3.a2s3_j.43$func$/openlane/designs/teras/src/arith_to_s3.v:95$95.$result[0] ));
 sky130_fd_sc_hd__or4_1 _10301_ (.A(\sa_inst._00_[0] ),
    .B(\sa_inst._00_[1] ),
    .C(\sa_inst._00_[7] ),
    .D(_00810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04319_));
 sky130_fd_sc_hd__clkbuf_1 _10302_ (.A(_04319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:2.a2s3_j._07_ ));
 sky130_fd_sc_hd__xnor2_1 _10303_ (.A(\sa_inst._00_[6] ),
    .B(\sa_inst._00_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_a2s3:2.a2s3_j.43$func$/openlane/designs/teras/src/arith_to_s3.v:95$95.$result[0] ));
 sky130_fd_sc_hd__xor2_1 _10304_ (.A(_02730_),
    .B(\sa_inst.sak._03_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04320_));
 sky130_fd_sc_hd__o21a_1 _10305_ (.A1(_02672_),
    .A2(\sa_inst.sak._03_[0] ),
    .B1(_04320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04321_));
 sky130_fd_sc_hd__nor3_1 _10306_ (.A(_02672_),
    .B(\sa_inst.sak._03_[0] ),
    .C(_04320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04322_));
 sky130_fd_sc_hd__nor2_1 _10307_ (.A(_04321_),
    .B(_04322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._08_[1] ));
 sky130_fd_sc_hd__a21oi_1 _10308_ (.A1(_02730_),
    .A2(\sa_inst.sak._03_[1] ),
    .B1(_04321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04323_));
 sky130_fd_sc_hd__nor2_1 _10309_ (.A(_02654_),
    .B(\sa_inst.sak._03_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04324_));
 sky130_fd_sc_hd__nand2_1 _10310_ (.A(_02654_),
    .B(\sa_inst.sak._03_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04325_));
 sky130_fd_sc_hd__and2b_1 _10311_ (.A_N(_04324_),
    .B(_04325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04326_));
 sky130_fd_sc_hd__xnor2_1 _10312_ (.A(_04323_),
    .B(_04326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._08_[2] ));
 sky130_fd_sc_hd__or2_1 _10313_ (.A(\sa_inst.sak._13_[3] ),
    .B(\sa_inst.sak._03_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04327_));
 sky130_fd_sc_hd__nand2_1 _10314_ (.A(\sa_inst.sak._13_[3] ),
    .B(\sa_inst.sak._03_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04328_));
 sky130_fd_sc_hd__nand2_1 _10315_ (.A(_04327_),
    .B(_04328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04329_));
 sky130_fd_sc_hd__o21ai_1 _10316_ (.A1(_04323_),
    .A2(_04324_),
    .B1(_04325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04330_));
 sky130_fd_sc_hd__xnor2_1 _10317_ (.A(_04329_),
    .B(_04330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._08_[3] ));
 sky130_fd_sc_hd__a21bo_1 _10318_ (.A1(_04327_),
    .A2(_04330_),
    .B1_N(_04328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._08_[4] ));
 sky130_fd_sc_hd__xnor2_1 _10319_ (.A(\sa_inst.cols_a2s3:3.a2s3_j._23_[1] ),
    .B(\sa_inst.sak._08_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04331_));
 sky130_fd_sc_hd__o21a_1 _10320_ (.A1(\sa_inst._07_[0] ),
    .A2(\sa_inst.sak._08_[0] ),
    .B1(_04331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04332_));
 sky130_fd_sc_hd__nor3_1 _10321_ (.A(\sa_inst._07_[0] ),
    .B(\sa_inst.sak._08_[0] ),
    .C(_04331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04333_));
 sky130_fd_sc_hd__nor2_1 _10322_ (.A(_04332_),
    .B(_04333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._08_[1] ));
 sky130_fd_sc_hd__a21oi_1 _10323_ (.A1(\sa_inst._07_[1] ),
    .A2(\sa_inst.sak._08_[1] ),
    .B1(_04332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04334_));
 sky130_fd_sc_hd__nor2_2 _10324_ (.A(\sa_inst.cols_a2s3:3.a2s3_j._23_[1] ),
    .B(\sa_inst.cols_a2s3:3.a2s3_j._23_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04335_));
 sky130_fd_sc_hd__and2_1 _10325_ (.A(\sa_inst.cols_a2s3:3.a2s3_j._23_[1] ),
    .B(\sa_inst.cols_a2s3:3.a2s3_j._23_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04336_));
 sky130_fd_sc_hd__or2_1 _10326_ (.A(_04335_),
    .B(_04336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04337_));
 sky130_fd_sc_hd__buf_2 _10327_ (.A(_04337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst._07_[2] ));
 sky130_fd_sc_hd__xor2_1 _10328_ (.A(\sa_inst.sak._08_[2] ),
    .B(\sa_inst._07_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04338_));
 sky130_fd_sc_hd__xnor2_1 _10329_ (.A(_04334_),
    .B(_04338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._08_[2] ));
 sky130_fd_sc_hd__xnor2_4 _10330_ (.A(\sa_inst.cols_a2s3:3.a2s3_j._23_[3] ),
    .B(_04335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst._07_[3] ));
 sky130_fd_sc_hd__xor2_1 _10331_ (.A(\sa_inst.sak._08_[3] ),
    .B(\sa_inst._07_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04339_));
 sky130_fd_sc_hd__a21bo_1 _10332_ (.A1(\sa_inst.sak._08_[2] ),
    .A2(\sa_inst._07_[2] ),
    .B1_N(_04334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04340_));
 sky130_fd_sc_hd__o21ai_1 _10333_ (.A1(\sa_inst.sak._08_[2] ),
    .A2(\sa_inst._07_[2] ),
    .B1(_04340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04341_));
 sky130_fd_sc_hd__xnor2_1 _10334_ (.A(_04339_),
    .B(_04341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._08_[3] ));
 sky130_fd_sc_hd__a21bo_1 _10335_ (.A1(\sa_inst.sak._08_[3] ),
    .A2(\sa_inst._07_[3] ),
    .B1_N(_04341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04342_));
 sky130_fd_sc_hd__o21a_1 _10336_ (.A1(\sa_inst.sak._08_[3] ),
    .A2(\sa_inst._07_[3] ),
    .B1(_04342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._08_[4] ));
 sky130_fd_sc_hd__xnor2_1 _10337_ (.A(\sa_inst.cols_a2s3:2.a2s3_j._23_[1] ),
    .B(_01199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04343_));
 sky130_fd_sc_hd__o21a_1 _10338_ (.A1(_01132_),
    .A2(\sa_inst._06_[0] ),
    .B1(_04343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04344_));
 sky130_fd_sc_hd__nor3_1 _10339_ (.A(_01132_),
    .B(\sa_inst._06_[0] ),
    .C(_04343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04345_));
 sky130_fd_sc_hd__nor2_1 _10340_ (.A(_04344_),
    .B(_04345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._08_[1] ));
 sky130_fd_sc_hd__a21oi_2 _10341_ (.A1(\sa_inst._06_[1] ),
    .A2(_01199_),
    .B1(_04344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04346_));
 sky130_fd_sc_hd__nor2_2 _10342_ (.A(\sa_inst.cols_a2s3:2.a2s3_j._23_[1] ),
    .B(\sa_inst.cols_a2s3:2.a2s3_j._23_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04347_));
 sky130_fd_sc_hd__and2_1 _10343_ (.A(\sa_inst.cols_a2s3:2.a2s3_j._23_[1] ),
    .B(\sa_inst.cols_a2s3:2.a2s3_j._23_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04348_));
 sky130_fd_sc_hd__or2_1 _10344_ (.A(_04347_),
    .B(_04348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04349_));
 sky130_fd_sc_hd__clkbuf_4 _10345_ (.A(_04349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst._06_[2] ));
 sky130_fd_sc_hd__xnor2_1 _10346_ (.A(_01060_),
    .B(\sa_inst._06_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04350_));
 sky130_fd_sc_hd__xnor2_1 _10347_ (.A(_04346_),
    .B(_04350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._08_[2] ));
 sky130_fd_sc_hd__xnor2_4 _10348_ (.A(\sa_inst.cols_a2s3:2.a2s3_j._23_[3] ),
    .B(_04347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst._06_[3] ));
 sky130_fd_sc_hd__xnor2_1 _10349_ (.A(_01072_),
    .B(\sa_inst._06_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04351_));
 sky130_fd_sc_hd__a21bo_1 _10350_ (.A1(_01144_),
    .A2(\sa_inst._06_[2] ),
    .B1_N(_04346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04352_));
 sky130_fd_sc_hd__o21ai_1 _10351_ (.A1(_01144_),
    .A2(\sa_inst._06_[2] ),
    .B1(_04352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04353_));
 sky130_fd_sc_hd__xnor2_1 _10352_ (.A(_04351_),
    .B(_04353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._08_[3] ));
 sky130_fd_sc_hd__a21bo_1 _10353_ (.A1(\sa_inst.sak._00_[3] ),
    .A2(\sa_inst._06_[3] ),
    .B1_N(_04353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04354_));
 sky130_fd_sc_hd__o21a_1 _10354_ (.A1(\sa_inst.sak._00_[3] ),
    .A2(\sa_inst._06_[3] ),
    .B1(_04354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._08_[4] ));
 sky130_fd_sc_hd__nor2_1 _10355_ (.A(\sa_inst.cols_a2s3:1.a2s3_j._23_[1] ),
    .B(\sa_inst.cols_a2s3:1.a2s3_j._23_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04355_));
 sky130_fd_sc_hd__and2_1 _10356_ (.A(\sa_inst.cols_a2s3:1.a2s3_j._23_[1] ),
    .B(\sa_inst.cols_a2s3:1.a2s3_j._23_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04356_));
 sky130_fd_sc_hd__or2_1 _10357_ (.A(_04355_),
    .B(_04356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04357_));
 sky130_fd_sc_hd__clkbuf_1 _10358_ (.A(_04357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst._05_[2] ));
 sky130_fd_sc_hd__xnor2_1 _10359_ (.A(\sa_inst.cols_a2s3:1.a2s3_j._23_[3] ),
    .B(_04355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst._05_[3] ));
 sky130_fd_sc_hd__clkbuf_1 _10360_ (.A(\sa_inst.sak._19_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04358_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10361_ (.A(\sa_inst.sak._19_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04359_));
 sky130_fd_sc_hd__clkbuf_1 _10362_ (.A(_04359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04360_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10363_ (.A(\sa_inst.sak._19_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04361_));
 sky130_fd_sc_hd__or2_1 _10364_ (.A(_04360_),
    .B(_04361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04362_));
 sky130_fd_sc_hd__nand2_1 _10365_ (.A(_04359_),
    .B(_04361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04363_));
 sky130_fd_sc_hd__and3_1 _10366_ (.A(_04358_),
    .B(_04362_),
    .C(_04363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04364_));
 sky130_fd_sc_hd__clkbuf_1 _10367_ (.A(_04364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w3_0 ));
 sky130_fd_sc_hd__inv_2 _10368_ (.A(\sa_inst.sak._19_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04365_));
 sky130_fd_sc_hd__clkbuf_2 _10369_ (.A(\sa_inst.sak._19_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04366_));
 sky130_fd_sc_hd__and2_1 _10370_ (.A(\sa_inst.sak._19_[4] ),
    .B(_04366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04367_));
 sky130_fd_sc_hd__nand3_1 _10371_ (.A(_04358_),
    .B(_04359_),
    .C(_04366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04368_));
 sky130_fd_sc_hd__o221a_1 _10372_ (.A1(_04358_),
    .A2(_04365_),
    .B1(_04367_),
    .B2(_04360_),
    .C1(_04368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w4_0 ));
 sky130_fd_sc_hd__clkbuf_1 _10373_ (.A(\sa_inst.sak._19_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04369_));
 sky130_fd_sc_hd__inv_2 _10374_ (.A(_04366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04370_));
 sky130_fd_sc_hd__o2bb2a_1 _10375_ (.A1_N(_04358_),
    .A2_N(_04369_),
    .B1(_04370_),
    .B2(_04365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04371_));
 sky130_fd_sc_hd__and3_1 _10376_ (.A(_04361_),
    .B(_04369_),
    .C(_04367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04372_));
 sky130_fd_sc_hd__nor2_1 _10377_ (.A(_04371_),
    .B(_04372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04373_));
 sky130_fd_sc_hd__and2_1 _10378_ (.A(_04363_),
    .B(_04368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04374_));
 sky130_fd_sc_hd__a21o_1 _10379_ (.A1(_04361_),
    .A2(_04367_),
    .B1(_04374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04375_));
 sky130_fd_sc_hd__xnor2_1 _10380_ (.A(_04373_),
    .B(_04375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w5_0 ));
 sky130_fd_sc_hd__a22o_1 _10381_ (.A1(\sa_inst.sak._19_[5] ),
    .A2(\sa_inst.sak._19_[8] ),
    .B1(\sa_inst.sak._19_[9] ),
    .B2(\sa_inst.sak._19_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04376_));
 sky130_fd_sc_hd__and4_1 _10382_ (.A(\sa_inst.sak._19_[4] ),
    .B(\sa_inst.sak._19_[5] ),
    .C(\sa_inst.sak._19_[8] ),
    .D(\sa_inst.sak._19_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04377_));
 sky130_fd_sc_hd__a31o_1 _10383_ (.A1(\sa_inst.sak._19_[6] ),
    .A2(\sa_inst.sak._19_[7] ),
    .A3(_04376_),
    .B1(_04377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04378_));
 sky130_fd_sc_hd__and2_1 _10384_ (.A(\sa_inst.sak._19_[7] ),
    .B(_04378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04379_));
 sky130_fd_sc_hd__o21ba_1 _10385_ (.A1(\sa_inst.sak._19_[7] ),
    .A2(_04377_),
    .B1_N(_04379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04380_));
 sky130_fd_sc_hd__nand2_1 _10386_ (.A(_04359_),
    .B(\sa_inst.sak._19_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04381_));
 sky130_fd_sc_hd__and2b_1 _10387_ (.A_N(_04377_),
    .B(_04376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04382_));
 sky130_fd_sc_hd__xnor2_1 _10388_ (.A(_04381_),
    .B(_04382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04383_));
 sky130_fd_sc_hd__and2_1 _10389_ (.A(_04380_),
    .B(_04383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04384_));
 sky130_fd_sc_hd__nor2_1 _10390_ (.A(_04380_),
    .B(_04383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04385_));
 sky130_fd_sc_hd__nor2_1 _10391_ (.A(_04384_),
    .B(_04385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04386_));
 sky130_fd_sc_hd__and2_1 _10392_ (.A(_04378_),
    .B(_04386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04387_));
 sky130_fd_sc_hd__nor2_1 _10393_ (.A(_04378_),
    .B(_04386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04388_));
 sky130_fd_sc_hd__nor2_1 _10394_ (.A(_04387_),
    .B(_04388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04389_));
 sky130_fd_sc_hd__and2_1 _10395_ (.A(_04372_),
    .B(_04389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04390_));
 sky130_fd_sc_hd__or2_1 _10396_ (.A(_04372_),
    .B(_04389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04391_));
 sky130_fd_sc_hd__or2b_1 _10397_ (.A(_04390_),
    .B_N(_04391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04392_));
 sky130_fd_sc_hd__and2b_1 _10398_ (.A_N(_04374_),
    .B(_04373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04393_));
 sky130_fd_sc_hd__a31o_1 _10399_ (.A1(_04360_),
    .A2(_04361_),
    .A3(_04366_),
    .B1(_04393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04394_));
 sky130_fd_sc_hd__xnor2_1 _10400_ (.A(_04392_),
    .B(_04394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w6_0 ));
 sky130_fd_sc_hd__clkbuf_1 _10401_ (.A(\sa_inst.sak._19_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04395_));
 sky130_fd_sc_hd__nand2_1 _10402_ (.A(_04369_),
    .B(_04395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04396_));
 sky130_fd_sc_hd__a22o_1 _10403_ (.A1(_04359_),
    .A2(\sa_inst.sak._19_[8] ),
    .B1(\sa_inst.sak._19_[9] ),
    .B2(\sa_inst.sak._19_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04397_));
 sky130_fd_sc_hd__o21a_1 _10404_ (.A1(_04363_),
    .A2(_04396_),
    .B1(_04397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04398_));
 sky130_fd_sc_hd__xnor2_1 _10405_ (.A(_04379_),
    .B(_04398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04399_));
 sky130_fd_sc_hd__o21ba_1 _10406_ (.A1(_04384_),
    .A2(_04387_),
    .B1_N(_04399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04400_));
 sky130_fd_sc_hd__or3b_1 _10407_ (.A(_04384_),
    .B(_04387_),
    .C_N(_04399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04401_));
 sky130_fd_sc_hd__and2b_1 _10408_ (.A_N(_04400_),
    .B(_04401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04402_));
 sky130_fd_sc_hd__a21oi_1 _10409_ (.A1(_04391_),
    .A2(_04394_),
    .B1(_04390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04403_));
 sky130_fd_sc_hd__xnor2_1 _10410_ (.A(_04402_),
    .B(_04403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w7_0 ));
 sky130_fd_sc_hd__and3_1 _10411_ (.A(_04389_),
    .B(_04393_),
    .C(_04401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04404_));
 sky130_fd_sc_hd__o2bb2a_1 _10412_ (.A1_N(_04379_),
    .A2_N(_04397_),
    .B1(_04396_),
    .B2(_04363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04405_));
 sky130_fd_sc_hd__and2_1 _10413_ (.A(_04369_),
    .B(_04370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04406_));
 sky130_fd_sc_hd__a21oi_1 _10414_ (.A1(_04360_),
    .A2(_04395_),
    .B1(_04406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04407_));
 sky130_fd_sc_hd__and3_1 _10415_ (.A(_04360_),
    .B(_04395_),
    .C(_04406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04408_));
 sky130_fd_sc_hd__nor2_1 _10416_ (.A(_04407_),
    .B(_04408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04409_));
 sky130_fd_sc_hd__and2b_1 _10417_ (.A_N(_04405_),
    .B(_04409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04410_));
 sky130_fd_sc_hd__and2b_1 _10418_ (.A_N(_04409_),
    .B(_04405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04411_));
 sky130_fd_sc_hd__nor2_1 _10419_ (.A(_04410_),
    .B(_04411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04412_));
 sky130_fd_sc_hd__o21a_1 _10420_ (.A1(_04400_),
    .A2(_04404_),
    .B1(_04412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04413_));
 sky130_fd_sc_hd__nor3_1 _10421_ (.A(_04400_),
    .B(_04404_),
    .C(_04412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04414_));
 sky130_fd_sc_hd__nor2_1 _10422_ (.A(_04413_),
    .B(_04414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w8_0 ));
 sky130_fd_sc_hd__or2_1 _10423_ (.A(_04369_),
    .B(_04395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04415_));
 sky130_fd_sc_hd__a31o_1 _10424_ (.A1(_04366_),
    .A2(_04396_),
    .A3(_04415_),
    .B1(_04408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04416_));
 sky130_fd_sc_hd__o21ai_1 _10425_ (.A1(_04410_),
    .A2(_04413_),
    .B1(_04416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04417_));
 sky130_fd_sc_hd__or3_1 _10426_ (.A(_04410_),
    .B(_04413_),
    .C(_04416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04418_));
 sky130_fd_sc_hd__and2_1 _10427_ (.A(_04417_),
    .B(_04418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04419_));
 sky130_fd_sc_hd__clkbuf_1 _10428_ (.A(_04419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w9_0 ));
 sky130_fd_sc_hd__and3b_1 _10429_ (.A_N(_04406_),
    .B(_04417_),
    .C(_04395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04420_));
 sky130_fd_sc_hd__clkbuf_1 _10430_ (.A(_04420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w10_0 ));
 sky130_fd_sc_hd__nand2_1 _10431_ (.A(_04396_),
    .B(_04417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w11_0 ));
 sky130_fd_sc_hd__nor2_1 _10432_ (.A(_04358_),
    .B(_04365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w2_0 ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10433_ (.A(\sa_inst.sak._07_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04421_));
 sky130_fd_sc_hd__clkbuf_2 _10434_ (.A(_04421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04422_));
 sky130_fd_sc_hd__inv_2 _10435_ (.A(_04422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04423_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10436_ (.A(\sa_inst.sak._07_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04424_));
 sky130_fd_sc_hd__inv_2 _10437_ (.A(\sa_inst.sak._07_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04425_));
 sky130_fd_sc_hd__nor2_1 _10438_ (.A(_04424_),
    .B(_04425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w2_0 ));
 sky130_fd_sc_hd__nor2_1 _10439_ (.A(_04423_),
    .B(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w2_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04426_));
 sky130_fd_sc_hd__clkbuf_2 _10440_ (.A(\sa_inst.sak._07_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04427_));
 sky130_fd_sc_hd__and2_1 _10441_ (.A(_04424_),
    .B(_04427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04428_));
 sky130_fd_sc_hd__mux2_1 _10442_ (.A0(_04426_),
    .A1(_04423_),
    .S(_04428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04429_));
 sky130_fd_sc_hd__clkbuf_1 _10443_ (.A(_04429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w4_0 ));
 sky130_fd_sc_hd__and3_1 _10444_ (.A(\sa_inst.sak._07_[5] ),
    .B(_04422_),
    .C(_04428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04430_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10445_ (.A(\sa_inst.sak._07_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04431_));
 sky130_fd_sc_hd__inv_2 _10446_ (.A(_04427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04432_));
 sky130_fd_sc_hd__o2bb2a_1 _10447_ (.A1_N(_04424_),
    .A2_N(_04431_),
    .B1(_04425_),
    .B2(_04432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04433_));
 sky130_fd_sc_hd__and2_1 _10448_ (.A(\sa_inst.sak._07_[8] ),
    .B(\sa_inst.sak._07_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04434_));
 sky130_fd_sc_hd__and2_1 _10449_ (.A(_04428_),
    .B(_04434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04435_));
 sky130_fd_sc_hd__or2_1 _10450_ (.A(_04433_),
    .B(_04435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04436_));
 sky130_fd_sc_hd__o21ai_1 _10451_ (.A1(\sa_inst.sak._07_[5] ),
    .A2(_04428_),
    .B1(_04422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04437_));
 sky130_fd_sc_hd__xnor2_1 _10452_ (.A(_04436_),
    .B(_04437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04438_));
 sky130_fd_sc_hd__xnor2_1 _10453_ (.A(_04430_),
    .B(_04438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w5_0 ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10454_ (.A(\sa_inst.sak._07_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04439_));
 sky130_fd_sc_hd__a21o_1 _10455_ (.A1(_04424_),
    .A2(_04439_),
    .B1(_04434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04440_));
 sky130_fd_sc_hd__and3_1 _10456_ (.A(\sa_inst.sak._07_[4] ),
    .B(\sa_inst.sak._07_[9] ),
    .C(_04434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04441_));
 sky130_fd_sc_hd__a31o_1 _10457_ (.A1(\sa_inst.sak._07_[7] ),
    .A2(\sa_inst.sak._07_[6] ),
    .A3(_04440_),
    .B1(_04441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04442_));
 sky130_fd_sc_hd__and2_1 _10458_ (.A(\sa_inst.sak._07_[7] ),
    .B(_04442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04443_));
 sky130_fd_sc_hd__o21ba_1 _10459_ (.A1(_04427_),
    .A2(_04441_),
    .B1_N(_04443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04444_));
 sky130_fd_sc_hd__nand2_1 _10460_ (.A(_04427_),
    .B(_04421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04445_));
 sky130_fd_sc_hd__and2b_1 _10461_ (.A_N(_04441_),
    .B(_04440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04446_));
 sky130_fd_sc_hd__xnor2_1 _10462_ (.A(_04445_),
    .B(_04446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04447_));
 sky130_fd_sc_hd__xor2_1 _10463_ (.A(_04444_),
    .B(_04447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04448_));
 sky130_fd_sc_hd__and2_1 _10464_ (.A(_04442_),
    .B(_04448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04449_));
 sky130_fd_sc_hd__nor2_1 _10465_ (.A(_04442_),
    .B(_04448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04450_));
 sky130_fd_sc_hd__nor2_1 _10466_ (.A(_04449_),
    .B(_04450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04451_));
 sky130_fd_sc_hd__and2_1 _10467_ (.A(_04435_),
    .B(_04451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04452_));
 sky130_fd_sc_hd__or2_1 _10468_ (.A(_04435_),
    .B(_04451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04453_));
 sky130_fd_sc_hd__or2b_1 _10469_ (.A(_04452_),
    .B_N(_04453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04454_));
 sky130_fd_sc_hd__o22ai_2 _10470_ (.A1(_04425_),
    .A2(_04445_),
    .B1(_04436_),
    .B2(_04437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04455_));
 sky130_fd_sc_hd__xnor2_1 _10471_ (.A(_04454_),
    .B(_04455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w6_0 ));
 sky130_fd_sc_hd__a21oi_1 _10472_ (.A1(_04444_),
    .A2(_04447_),
    .B1(_04449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04456_));
 sky130_fd_sc_hd__a22o_1 _10473_ (.A1(_04431_),
    .A2(_04421_),
    .B1(_04439_),
    .B2(\sa_inst.sak._07_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04457_));
 sky130_fd_sc_hd__inv_2 _10474_ (.A(_04457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04458_));
 sky130_fd_sc_hd__a31o_1 _10475_ (.A1(_04421_),
    .A2(_04439_),
    .A3(_04434_),
    .B1(_04458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04459_));
 sky130_fd_sc_hd__xor2_1 _10476_ (.A(_04443_),
    .B(_04459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04460_));
 sky130_fd_sc_hd__xnor2_1 _10477_ (.A(_04456_),
    .B(_04460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04461_));
 sky130_fd_sc_hd__a21oi_1 _10478_ (.A1(_04453_),
    .A2(_04455_),
    .B1(_04452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04462_));
 sky130_fd_sc_hd__xor2_1 _10479_ (.A(_04461_),
    .B(_04462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w7_0 ));
 sky130_fd_sc_hd__nor2_1 _10480_ (.A(_04456_),
    .B(_04460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04463_));
 sky130_fd_sc_hd__nor2_1 _10481_ (.A(_04461_),
    .B(_04462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04464_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10482_ (.A(_04439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04465_));
 sky130_fd_sc_hd__and2_1 _10483_ (.A(_04431_),
    .B(_04432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04466_));
 sky130_fd_sc_hd__a21oi_1 _10484_ (.A1(_04422_),
    .A2(_04465_),
    .B1(_04466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04467_));
 sky130_fd_sc_hd__and3_1 _10485_ (.A(_04421_),
    .B(_04439_),
    .C(_04466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04468_));
 sky130_fd_sc_hd__or2_1 _10486_ (.A(_04467_),
    .B(_04468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04469_));
 sky130_fd_sc_hd__a32o_1 _10487_ (.A1(_04422_),
    .A2(_04465_),
    .A3(_04434_),
    .B1(_04443_),
    .B2(_04457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04470_));
 sky130_fd_sc_hd__xnor2_1 _10488_ (.A(_04469_),
    .B(_04470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04471_));
 sky130_fd_sc_hd__o21ai_1 _10489_ (.A1(_04463_),
    .A2(_04464_),
    .B1(_04471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04472_));
 sky130_fd_sc_hd__or3_1 _10490_ (.A(_04463_),
    .B(_04464_),
    .C(_04471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04473_));
 sky130_fd_sc_hd__and2_1 _10491_ (.A(_04472_),
    .B(_04473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04474_));
 sky130_fd_sc_hd__clkbuf_1 _10492_ (.A(_04474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w8_0 ));
 sky130_fd_sc_hd__or2b_1 _10493_ (.A(_04469_),
    .B_N(_04470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04475_));
 sky130_fd_sc_hd__or2_1 _10494_ (.A(_04431_),
    .B(_04465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04476_));
 sky130_fd_sc_hd__nand2_1 _10495_ (.A(_04431_),
    .B(_04465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04477_));
 sky130_fd_sc_hd__a31oi_1 _10496_ (.A1(_04427_),
    .A2(_04476_),
    .A3(_04477_),
    .B1(_04468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04478_));
 sky130_fd_sc_hd__a21o_1 _10497_ (.A1(_04475_),
    .A2(_04472_),
    .B1(_04478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04479_));
 sky130_fd_sc_hd__nand3_1 _10498_ (.A(_04475_),
    .B(_04472_),
    .C(_04478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04480_));
 sky130_fd_sc_hd__and2_1 _10499_ (.A(_04479_),
    .B(_04480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04481_));
 sky130_fd_sc_hd__clkbuf_1 _10500_ (.A(_04481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w9_0 ));
 sky130_fd_sc_hd__and3b_1 _10501_ (.A_N(_04466_),
    .B(_04479_),
    .C(_04465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04482_));
 sky130_fd_sc_hd__clkbuf_1 _10502_ (.A(_04482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w10_0 ));
 sky130_fd_sc_hd__nand2_1 _10503_ (.A(_04477_),
    .B(_04479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w11_0 ));
 sky130_fd_sc_hd__o21ai_1 _10504_ (.A1(_04425_),
    .A2(_04423_),
    .B1(_04424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04483_));
 sky130_fd_sc_hd__a21oi_1 _10505_ (.A1(_04425_),
    .A2(_04423_),
    .B1(_04483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w3_0 ));
 sky130_fd_sc_hd__inv_2 _10506_ (.A(\sa_inst._05_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04484_));
 sky130_fd_sc_hd__clkbuf_1 _10507_ (.A(\sa_inst._05_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04485_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10508_ (.A(\sa_inst._05_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04486_));
 sky130_fd_sc_hd__inv_2 _10509_ (.A(_04486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04487_));
 sky130_fd_sc_hd__nor2_1 _10510_ (.A(_04485_),
    .B(_04487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w2_0 ));
 sky130_fd_sc_hd__nor2_1 _10511_ (.A(_04484_),
    .B(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w2_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04488_));
 sky130_fd_sc_hd__and2_1 _10512_ (.A(_04485_),
    .B(\sa_inst._05_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04489_));
 sky130_fd_sc_hd__mux2_1 _10513_ (.A0(_04488_),
    .A1(_04484_),
    .S(_04489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04490_));
 sky130_fd_sc_hd__clkbuf_1 _10514_ (.A(_04490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w4_0 ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10515_ (.A(\sa_inst._05_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04491_));
 sky130_fd_sc_hd__inv_2 _10516_ (.A(\sa_inst._05_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04492_));
 sky130_fd_sc_hd__o2bb2a_1 _10517_ (.A1_N(_04485_),
    .A2_N(_04491_),
    .B1(_04487_),
    .B2(_04492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04493_));
 sky130_fd_sc_hd__and2_1 _10518_ (.A(\sa_inst._05_[8] ),
    .B(\sa_inst._05_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04494_));
 sky130_fd_sc_hd__and2_1 _10519_ (.A(_04489_),
    .B(_04494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04495_));
 sky130_fd_sc_hd__or2_1 _10520_ (.A(_04493_),
    .B(_04495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04496_));
 sky130_fd_sc_hd__nor2_1 _10521_ (.A(_04492_),
    .B(_04484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04497_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10522_ (.A(\sa_inst._05_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04498_));
 sky130_fd_sc_hd__o21ai_1 _10523_ (.A1(_04486_),
    .A2(_04489_),
    .B1(_04498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04499_));
 sky130_fd_sc_hd__a31o_1 _10524_ (.A1(_04485_),
    .A2(_04486_),
    .A3(_04497_),
    .B1(_04499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04500_));
 sky130_fd_sc_hd__xor2_1 _10525_ (.A(_04496_),
    .B(_04500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w5_0 ));
 sky130_fd_sc_hd__and3_1 _10526_ (.A(\sa_inst._05_[4] ),
    .B(\sa_inst._05_[9] ),
    .C(_04494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04501_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10527_ (.A(\sa_inst._05_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04502_));
 sky130_fd_sc_hd__a21o_1 _10528_ (.A1(\sa_inst._05_[4] ),
    .A2(_04502_),
    .B1(_04494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04503_));
 sky130_fd_sc_hd__o21a_1 _10529_ (.A1(_04497_),
    .A2(_04501_),
    .B1(_04503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04504_));
 sky130_fd_sc_hd__and2_1 _10530_ (.A(\sa_inst._05_[7] ),
    .B(_04504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04505_));
 sky130_fd_sc_hd__nor2_1 _10531_ (.A(\sa_inst._05_[7] ),
    .B(_04501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04506_));
 sky130_fd_sc_hd__and2b_1 _10532_ (.A_N(_04501_),
    .B(_04503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04507_));
 sky130_fd_sc_hd__xor2_1 _10533_ (.A(_04497_),
    .B(_04507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04508_));
 sky130_fd_sc_hd__or3b_1 _10534_ (.A(_04505_),
    .B(_04506_),
    .C_N(_04508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04509_));
 sky130_fd_sc_hd__o21bai_1 _10535_ (.A1(_04505_),
    .A2(_04506_),
    .B1_N(_04508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04510_));
 sky130_fd_sc_hd__nand2_1 _10536_ (.A(_04509_),
    .B(_04510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04511_));
 sky130_fd_sc_hd__xnor2_1 _10537_ (.A(_04504_),
    .B(_04511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04512_));
 sky130_fd_sc_hd__and2_1 _10538_ (.A(_04495_),
    .B(_04512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04513_));
 sky130_fd_sc_hd__or2_1 _10539_ (.A(_04495_),
    .B(_04512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04514_));
 sky130_fd_sc_hd__or2b_1 _10540_ (.A(_04513_),
    .B_N(_04514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04515_));
 sky130_fd_sc_hd__a2bb2o_1 _10541_ (.A1_N(_04496_),
    .A2_N(_04499_),
    .B1(_04497_),
    .B2(_04486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04516_));
 sky130_fd_sc_hd__xnor2_1 _10542_ (.A(_04515_),
    .B(_04516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w6_0 ));
 sky130_fd_sc_hd__o21ai_1 _10543_ (.A1(_04492_),
    .A2(_04498_),
    .B1(_04501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04517_));
 sky130_fd_sc_hd__a22o_1 _10544_ (.A1(_04491_),
    .A2(\sa_inst._05_[6] ),
    .B1(_04502_),
    .B2(_04486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04518_));
 sky130_fd_sc_hd__inv_2 _10545_ (.A(_04518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04519_));
 sky130_fd_sc_hd__a31o_1 _10546_ (.A1(\sa_inst._05_[6] ),
    .A2(_04502_),
    .A3(_04494_),
    .B1(_04519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04520_));
 sky130_fd_sc_hd__xor2_1 _10547_ (.A(_04505_),
    .B(_04520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04521_));
 sky130_fd_sc_hd__a21oi_1 _10548_ (.A1(_04509_),
    .A2(_04517_),
    .B1(_04521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04522_));
 sky130_fd_sc_hd__and3_1 _10549_ (.A(_04509_),
    .B(_04517_),
    .C(_04521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04523_));
 sky130_fd_sc_hd__or2_1 _10550_ (.A(_04522_),
    .B(_04523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04524_));
 sky130_fd_sc_hd__a21oi_1 _10551_ (.A1(_04514_),
    .A2(_04516_),
    .B1(_04513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04525_));
 sky130_fd_sc_hd__xor2_1 _10552_ (.A(_04524_),
    .B(_04525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w7_0 ));
 sky130_fd_sc_hd__nor2_1 _10553_ (.A(_04524_),
    .B(_04525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04526_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10554_ (.A(_04502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04527_));
 sky130_fd_sc_hd__and2_1 _10555_ (.A(_04491_),
    .B(_04492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04528_));
 sky130_fd_sc_hd__a21oi_1 _10556_ (.A1(_04498_),
    .A2(_04527_),
    .B1(_04528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04529_));
 sky130_fd_sc_hd__and3_1 _10557_ (.A(_04498_),
    .B(_04502_),
    .C(_04528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04530_));
 sky130_fd_sc_hd__or2_1 _10558_ (.A(_04529_),
    .B(_04530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04531_));
 sky130_fd_sc_hd__a32o_1 _10559_ (.A1(_04498_),
    .A2(_04527_),
    .A3(_04494_),
    .B1(_04505_),
    .B2(_04518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04532_));
 sky130_fd_sc_hd__xnor2_1 _10560_ (.A(_04531_),
    .B(_04532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04533_));
 sky130_fd_sc_hd__o21ai_1 _10561_ (.A1(_04522_),
    .A2(_04526_),
    .B1(_04533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04534_));
 sky130_fd_sc_hd__or3_1 _10562_ (.A(_04522_),
    .B(_04526_),
    .C(_04533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04535_));
 sky130_fd_sc_hd__and2_1 _10563_ (.A(_04534_),
    .B(_04535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04536_));
 sky130_fd_sc_hd__clkbuf_1 _10564_ (.A(_04536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w8_0 ));
 sky130_fd_sc_hd__or2b_1 _10565_ (.A(_04531_),
    .B_N(_04532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04537_));
 sky130_fd_sc_hd__or2_1 _10566_ (.A(_04491_),
    .B(_04527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04538_));
 sky130_fd_sc_hd__nand2_1 _10567_ (.A(_04491_),
    .B(_04527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04539_));
 sky130_fd_sc_hd__a31oi_1 _10568_ (.A1(\sa_inst._05_[7] ),
    .A2(_04538_),
    .A3(_04539_),
    .B1(_04530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04540_));
 sky130_fd_sc_hd__a21o_1 _10569_ (.A1(_04537_),
    .A2(_04534_),
    .B1(_04540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04541_));
 sky130_fd_sc_hd__nand3_1 _10570_ (.A(_04537_),
    .B(_04534_),
    .C(_04540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04542_));
 sky130_fd_sc_hd__and2_1 _10571_ (.A(_04541_),
    .B(_04542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04543_));
 sky130_fd_sc_hd__clkbuf_1 _10572_ (.A(_04543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w9_0 ));
 sky130_fd_sc_hd__and3b_1 _10573_ (.A_N(_04528_),
    .B(_04541_),
    .C(_04527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04544_));
 sky130_fd_sc_hd__clkbuf_1 _10574_ (.A(_04544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w10_0 ));
 sky130_fd_sc_hd__nand2_1 _10575_ (.A(_04539_),
    .B(_04541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w11_0 ));
 sky130_fd_sc_hd__o21ai_1 _10576_ (.A1(_04487_),
    .A2(_04484_),
    .B1(_04485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04545_));
 sky130_fd_sc_hd__a21oi_1 _10577_ (.A1(_04487_),
    .A2(_04484_),
    .B1(_04545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w3_0 ));
 sky130_fd_sc_hd__o31a_1 _10578_ (.A1(\sa_inst.sak._00_[11] ),
    .A2(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._25_ ),
    .A3(\sa_inst.sak.rows:1.cols:1.pe_ij._02_ ),
    .B1(_01198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._20_ ));
 sky130_fd_sc_hd__or2_1 _10579_ (.A(\sa_inst.sak._00_[11] ),
    .B(\sa_inst._06_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04546_));
 sky130_fd_sc_hd__clkbuf_1 _10580_ (.A(_04546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._02_ ));
 sky130_fd_sc_hd__o31a_1 _10581_ (.A1(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._11_ ),
    .A2(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._25_ ),
    .A3(\sa_inst.sak.rows:1.cols:2.pe_ij._02_ ),
    .B1(_01494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._20_ ));
 sky130_fd_sc_hd__or2_1 _10582_ (.A(\sa_inst._07_[11] ),
    .B(\sa_inst.sak._08_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04547_));
 sky130_fd_sc_hd__clkbuf_1 _10583_ (.A(_04547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._02_ ));
 sky130_fd_sc_hd__o31a_1 _10584_ (.A1(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._11_ ),
    .A2(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._25_ ),
    .A3(\sa_inst.sak.rows:1.cols:3.pe_ij._02_ ),
    .B1(_01927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._20_ ));
 sky130_fd_sc_hd__o31a_1 _10585_ (.A1(\sa_inst.sak.rows:2.cols:1.pe_ij._02_ ),
    .A2(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._11_ ),
    .A3(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._25_ ),
    .B1(_01494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._20_ ));
 sky130_fd_sc_hd__o31a_1 _10586_ (.A1(\sa_inst.sak.rows:2.cols:2.pe_ij._02_ ),
    .A2(\sa_inst.sak._13_[11] ),
    .A3(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._25_ ),
    .B1(_01927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._20_ ));
 sky130_fd_sc_hd__or2_1 _10587_ (.A(\sa_inst.sak._13_[11] ),
    .B(\sa_inst.sak._03_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04548_));
 sky130_fd_sc_hd__clkbuf_1 _10588_ (.A(_04548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._02_ ));
 sky130_fd_sc_hd__o31a_1 _10589_ (.A1(\sa_inst.sak.rows:2.cols:3.pe_ij._02_ ),
    .A2(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._11_ ),
    .A3(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._25_ ),
    .B1(_02878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._20_ ));
 sky130_fd_sc_hd__o31a_1 _10590_ (.A1(\sa_inst.sak.rows:3.cols:1.pe_ij._02_ ),
    .A2(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._11_ ),
    .A3(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._25_ ),
    .B1(_01927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._20_ ));
 sky130_fd_sc_hd__o31a_1 _10591_ (.A1(\sa_inst.sak.rows:3.cols:2.pe_ij._02_ ),
    .A2(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._11_ ),
    .A3(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._25_ ),
    .B1(_02878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._20_ ));
 sky130_fd_sc_hd__xor2_1 _10592_ (.A(\sa_inst.cols_a2s3:3.a2s3_j._15_[3] ),
    .B(_04307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:3.a2s3_j._15_[0] ));
 sky130_fd_sc_hd__xor2_1 _10593_ (.A(_04302_),
    .B(\sa_inst.cols_a2s3:3.a2s3_j._15_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:3.a2s3_j._15_[1] ));
 sky130_fd_sc_hd__xor2_1 _10594_ (.A(\sa_inst.cols_a2s3:3.a2s3_j._15_[3] ),
    .B(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._08_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:3.a2s3_j._15_[2] ));
 sky130_fd_sc_hd__o31a_1 _10595_ (.A1(\sa_inst.sak.rows:3.cols:3.pe_ij._02_ ),
    .A2(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._11_ ),
    .A3(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._25_ ),
    .B1(_03976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._20_ ));
 sky130_fd_sc_hd__xor2_1 _10596_ (.A(\sa_inst.cols_a2s3:2.a2s3_j._15_[3] ),
    .B(_04125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:2.a2s3_j._15_[0] ));
 sky130_fd_sc_hd__xor2_1 _10597_ (.A(_04120_),
    .B(\sa_inst.cols_a2s3:2.a2s3_j._15_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:2.a2s3_j._15_[1] ));
 sky130_fd_sc_hd__xor2_1 _10598_ (.A(\sa_inst.cols_a2s3:2.a2s3_j._15_[3] ),
    .B(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._08_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:2.a2s3_j._15_[2] ));
 sky130_fd_sc_hd__or4b_1 _10599_ (.A(\sa_inst._00_[0] ),
    .B(_00810_),
    .C(\sa_inst._00_[1] ),
    .D_N(\sa_inst._00_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04549_));
 sky130_fd_sc_hd__inv_2 _10600_ (.A(_04549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_a2s3:2.a2s3_j._05_ ));
 sky130_fd_sc_hd__and3_1 _10601_ (.A(_00817_),
    .B(\sa_inst.arith_in_col_0[7] ),
    .C(_04316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04550_));
 sky130_fd_sc_hd__clkbuf_1 _10602_ (.A(_04550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:1.a2s3_j._05_ ));
 sky130_fd_sc_hd__and2_1 _10603_ (.A(\sa_inst.cols_l2a:3.l2a_i.rshift._11_[0] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.rshift._18_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04551_));
 sky130_fd_sc_hd__or4_1 _10604_ (.A(\sa_inst.cols_l2a:3.l2a_i.rshift._27_ ),
    .B(\sa_inst.cols_l2a:3.l2a_i._04_[0] ),
    .C(\sa_inst.cols_l2a:3.l2a_i._01_ ),
    .D(\sa_inst.cols_l2a:3.l2a_i._08_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04552_));
 sky130_fd_sc_hd__o21a_1 _10605_ (.A1(_04551_),
    .A2(_04552_),
    .B1(\sa_inst.cols_l2a:3.l2a_i._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._46_ ));
 sky130_fd_sc_hd__or4_1 _10606_ (.A(_00849_),
    .B(_00852_),
    .C(_04151_),
    .D(_04156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04553_));
 sky130_fd_sc_hd__or3_1 _10607_ (.A(_04152_),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[16] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._08_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04554_));
 sky130_fd_sc_hd__or3b_1 _10608_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._09_ ),
    .B(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[8] ),
    .C_N(_04152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04555_));
 sky130_fd_sc_hd__a221o_1 _10609_ (.A1(_04154_),
    .A2(_04553_),
    .B1(_04554_),
    .B2(_04555_),
    .C1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._67_ ));
 sky130_fd_sc_hd__or4_1 _10610_ (.A(\sa_inst.cols_l2a:3.l2a_i.rshift._25_[1] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.rshift._25_[0] ),
    .C(\sa_inst.cols_l2a:3.l2a_i.rshift._25_[3] ),
    .D(\sa_inst.cols_l2a:3.l2a_i.rshift._25_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04556_));
 sky130_fd_sc_hd__or2_1 _10611_ (.A(\sa_inst.cols_l2a:3.l2a_i.rshift._26_[1] ),
    .B(\sa_inst.cols_l2a:3.l2a_i.rshift._26_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04557_));
 sky130_fd_sc_hd__a221o_1 _10612_ (.A1(\sa_inst.cols_l2a:3.l2a_i.rshift._00_[2] ),
    .A2(_04556_),
    .B1(_04557_),
    .B2(\sa_inst.cols_l2a:3.l2a_i.rshift._00_[1] ),
    .C1(\sa_inst.cols_l2a:3.l2a_i.rshift._22_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i.rshift._14_ ));
 sky130_fd_sc_hd__and2_1 _10613_ (.A(\sa_inst.cols_l2a:2.l2a_i.rshift._11_[0] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.rshift._18_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04558_));
 sky130_fd_sc_hd__or4_1 _10614_ (.A(\sa_inst.cols_l2a:2.l2a_i.rshift._27_ ),
    .B(\sa_inst.cols_l2a:2.l2a_i._04_[0] ),
    .C(\sa_inst.cols_l2a:2.l2a_i._01_ ),
    .D(\sa_inst.cols_l2a:2.l2a_i._08_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04559_));
 sky130_fd_sc_hd__o21a_1 _10615_ (.A1(_04558_),
    .A2(_04559_),
    .B1(\sa_inst.cols_l2a:2.l2a_i._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._46_ ));
 sky130_fd_sc_hd__or4_1 _10616_ (.A(_00899_),
    .B(_00902_),
    .C(_04203_),
    .D(_04208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04560_));
 sky130_fd_sc_hd__or3_1 _10617_ (.A(_04204_),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[16] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._08_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04561_));
 sky130_fd_sc_hd__or3b_1 _10618_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._09_ ),
    .B(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[8] ),
    .C_N(_04204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04562_));
 sky130_fd_sc_hd__a221o_1 _10619_ (.A1(_04206_),
    .A2(_04560_),
    .B1(_04561_),
    .B2(_04562_),
    .C1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._67_ ));
 sky130_fd_sc_hd__or4_1 _10620_ (.A(\sa_inst.cols_l2a:2.l2a_i.rshift._25_[1] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.rshift._25_[0] ),
    .C(\sa_inst.cols_l2a:2.l2a_i.rshift._25_[3] ),
    .D(\sa_inst.cols_l2a:2.l2a_i.rshift._25_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04563_));
 sky130_fd_sc_hd__or2_1 _10621_ (.A(\sa_inst.cols_l2a:2.l2a_i.rshift._26_[1] ),
    .B(\sa_inst.cols_l2a:2.l2a_i.rshift._26_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04564_));
 sky130_fd_sc_hd__a221o_1 _10622_ (.A1(\sa_inst.cols_l2a:2.l2a_i.rshift._00_[2] ),
    .A2(_04563_),
    .B1(_04564_),
    .B2(\sa_inst.cols_l2a:2.l2a_i.rshift._00_[1] ),
    .C1(\sa_inst.cols_l2a:2.l2a_i.rshift._22_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i.rshift._14_ ));
 sky130_fd_sc_hd__and2_1 _10623_ (.A(\sa_inst.cols_l2a:1.l2a_i.rshift._11_[0] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.rshift._18_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04565_));
 sky130_fd_sc_hd__or4_1 _10624_ (.A(\sa_inst.cols_l2a:1.l2a_i.rshift._27_ ),
    .B(\sa_inst.cols_l2a:1.l2a_i._04_[0] ),
    .C(\sa_inst.cols_l2a:1.l2a_i._01_ ),
    .D(\sa_inst.cols_l2a:1.l2a_i._08_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04566_));
 sky130_fd_sc_hd__o21a_1 _10625_ (.A1(_04565_),
    .A2(_04566_),
    .B1(\sa_inst.cols_l2a:1.l2a_i._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._46_ ));
 sky130_fd_sc_hd__or4_1 _10626_ (.A(_00949_),
    .B(_00952_),
    .C(_04255_),
    .D(_04260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04567_));
 sky130_fd_sc_hd__or3_1 _10627_ (.A(_04256_),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[16] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._08_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04568_));
 sky130_fd_sc_hd__or3b_1 _10628_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._09_ ),
    .B(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[8] ),
    .C_N(_04256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04569_));
 sky130_fd_sc_hd__a221o_1 _10629_ (.A1(_04258_),
    .A2(_04567_),
    .B1(_04568_),
    .B2(_04569_),
    .C1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._67_ ));
 sky130_fd_sc_hd__or4_1 _10630_ (.A(\sa_inst.cols_l2a:1.l2a_i.rshift._25_[1] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.rshift._25_[0] ),
    .C(\sa_inst.cols_l2a:1.l2a_i.rshift._25_[3] ),
    .D(\sa_inst.cols_l2a:1.l2a_i.rshift._25_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04570_));
 sky130_fd_sc_hd__or2_1 _10631_ (.A(\sa_inst.cols_l2a:1.l2a_i.rshift._26_[1] ),
    .B(\sa_inst.cols_l2a:1.l2a_i.rshift._26_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04571_));
 sky130_fd_sc_hd__a221o_1 _10632_ (.A1(\sa_inst.cols_l2a:1.l2a_i.rshift._00_[2] ),
    .A2(_04570_),
    .B1(_04571_),
    .B2(\sa_inst.cols_l2a:1.l2a_i.rshift._00_[1] ),
    .C1(\sa_inst.cols_l2a:1.l2a_i.rshift._22_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i.rshift._14_ ));
 sky130_fd_sc_hd__or4b_1 _10633_ (.A(\sa_inst._17_[0] ),
    .B(_00806_),
    .C(\sa_inst._17_[1] ),
    .D_N(\sa_inst._17_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04572_));
 sky130_fd_sc_hd__clkinv_2 _10634_ (.A(_04572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_a2s3:3.a2s3_j._05_ ));
 sky130_fd_sc_hd__xor2_1 _10635_ (.A(\sa_inst.cols_a2s3:1.a2s3_j._15_[3] ),
    .B(_04138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:1.a2s3_j._15_[0] ));
 sky130_fd_sc_hd__xor2_1 _10636_ (.A(_04133_),
    .B(\sa_inst.cols_a2s3:1.a2s3_j._15_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:1.a2s3_j._15_[1] ));
 sky130_fd_sc_hd__xor2_1 _10637_ (.A(\sa_inst.cols_a2s3:1.a2s3_j._15_[3] ),
    .B(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._08_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_a2s3:1.a2s3_j._15_[2] ));
 sky130_fd_sc_hd__xor2_1 _10638_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._07_ ),
    .B(\sa_inst.cols_l2a:3.l2a_i._31_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:3.l2a_i._31_[3] ));
 sky130_fd_sc_hd__o21ai_1 _10639_ (.A1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._07_ ),
    .A2(\sa_inst.cols_l2a:3.l2a_i._31_[2] ),
    .B1(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._01_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04573_));
 sky130_fd_sc_hd__xnor2_1 _10640_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._55_ ),
    .B(_04573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:3.l2a_i._31_[5] ));
 sky130_fd_sc_hd__xor2_1 _10641_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._07_ ),
    .B(\sa_inst.cols_l2a:2.l2a_i._31_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:2.l2a_i._31_[3] ));
 sky130_fd_sc_hd__o21ai_1 _10642_ (.A1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._07_ ),
    .A2(\sa_inst.cols_l2a:2.l2a_i._31_[2] ),
    .B1(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._01_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04574_));
 sky130_fd_sc_hd__xnor2_1 _10643_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._55_ ),
    .B(_04574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:2.l2a_i._31_[5] ));
 sky130_fd_sc_hd__xor2_1 _10644_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._07_ ),
    .B(\sa_inst.cols_l2a:1.l2a_i._31_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\sa_inst.cols_l2a:1.l2a_i._31_[3] ));
 sky130_fd_sc_hd__o21ai_1 _10645_ (.A1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._07_ ),
    .A2(\sa_inst.cols_l2a:1.l2a_i._31_[2] ),
    .B1(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._01_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04575_));
 sky130_fd_sc_hd__xnor2_1 _10646_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._55_ ),
    .B(_04575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\sa_inst.cols_l2a:1.l2a_i._31_[5] ));
 sky130_fd_sc_hd__and2_1 _10647_ (.A(_01626_),
    .B(_01617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04576_));
 sky130_fd_sc_hd__clkbuf_1 _10648_ (.A(_04576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00000_));
 sky130_fd_sc_hd__and2_1 _10649_ (.A(\sa_inst._12_[0] ),
    .B(_00802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04577_));
 sky130_fd_sc_hd__clkbuf_1 _10650_ (.A(_04577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00001_));
 sky130_fd_sc_hd__and2_1 _10651_ (.A(\sa_inst._12_[33] ),
    .B(_00762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04578_));
 sky130_fd_sc_hd__clkbuf_1 _10652_ (.A(_04578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00002_));
 sky130_fd_sc_hd__and2_1 _10653_ (.A(\sa_inst._12_[66] ),
    .B(_00722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04579_));
 sky130_fd_sc_hd__clkbuf_1 _10654_ (.A(_04579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00003_));
 sky130_fd_sc_hd__nor2_1 _10655_ (.A(\sa_inst.cols_l2a:1.l2a_i._27_ ),
    .B(\sa_inst.cols_l2a:1.l2a_i._23_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04580_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10656_ (.A(_04580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04581_));
 sky130_fd_sc_hd__o21ai_1 _10657_ (.A1(\sa_inst.cols_l2a:1.l2a_i._09_[0] ),
    .A2(\sa_inst.cols_l2a:1.l2a_i._15_ ),
    .B1(_04581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04582_));
 sky130_fd_sc_hd__a21oi_2 _10658_ (.A1(\sa_inst.cols_l2a:1.l2a_i._09_[0] ),
    .A2(\sa_inst.cols_l2a:1.l2a_i._15_ ),
    .B1(_04582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00004_));
 sky130_fd_sc_hd__and3_1 _10659_ (.A(\sa_inst.cols_l2a:1.l2a_i._09_[0] ),
    .B(\sa_inst.cols_l2a:1.l2a_i._15_ ),
    .C(\sa_inst.cols_l2a:1.l2a_i._09_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04583_));
 sky130_fd_sc_hd__a21o_1 _10660_ (.A1(\sa_inst.cols_l2a:1.l2a_i._09_[0] ),
    .A2(\sa_inst.cols_l2a:1.l2a_i._15_ ),
    .B1(\sa_inst.cols_l2a:1.l2a_i._09_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04584_));
 sky130_fd_sc_hd__and3b_1 _10661_ (.A_N(_04583_),
    .B(_04580_),
    .C(_04584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04585_));
 sky130_fd_sc_hd__clkbuf_1 _10662_ (.A(_04585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00005_));
 sky130_fd_sc_hd__and2_1 _10663_ (.A(\sa_inst.cols_l2a:1.l2a_i._09_[2] ),
    .B(_04583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04586_));
 sky130_fd_sc_hd__o21ai_1 _10664_ (.A1(\sa_inst.cols_l2a:1.l2a_i._09_[2] ),
    .A2(_04583_),
    .B1(_04581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04587_));
 sky130_fd_sc_hd__nor2_1 _10665_ (.A(_04586_),
    .B(_04587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00006_));
 sky130_fd_sc_hd__and3_1 _10666_ (.A(\sa_inst.cols_l2a:1.l2a_i._09_[2] ),
    .B(\sa_inst.cols_l2a:1.l2a_i._09_[3] ),
    .C(_04583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04588_));
 sky130_fd_sc_hd__o21ai_1 _10667_ (.A1(\sa_inst.cols_l2a:1.l2a_i._09_[3] ),
    .A2(_04586_),
    .B1(_04581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04589_));
 sky130_fd_sc_hd__nor2_1 _10668_ (.A(_04588_),
    .B(_04589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00007_));
 sky130_fd_sc_hd__o21ai_1 _10669_ (.A1(\sa_inst.cols_l2a:1.l2a_i._09_[4] ),
    .A2(_04588_),
    .B1(_04581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04590_));
 sky130_fd_sc_hd__a21oi_1 _10670_ (.A1(\sa_inst.cols_l2a:1.l2a_i._09_[4] ),
    .A2(_04588_),
    .B1(_04590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00008_));
 sky130_fd_sc_hd__and3_1 _10671_ (.A(\sa_inst.cols_l2a:1.l2a_i._09_[4] ),
    .B(\sa_inst.cols_l2a:1.l2a_i._09_[5] ),
    .C(_04588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04591_));
 sky130_fd_sc_hd__a21o_1 _10672_ (.A1(\sa_inst.cols_l2a:1.l2a_i._09_[4] ),
    .A2(_04588_),
    .B1(\sa_inst.cols_l2a:1.l2a_i._09_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04592_));
 sky130_fd_sc_hd__and3b_1 _10673_ (.A_N(_04591_),
    .B(_04580_),
    .C(_04592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04593_));
 sky130_fd_sc_hd__clkbuf_1 _10674_ (.A(_04593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00009_));
 sky130_fd_sc_hd__a21boi_1 _10675_ (.A1(\sa_inst.cols_l2a:1.l2a_i._09_[6] ),
    .A2(_04591_),
    .B1_N(_04581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04594_));
 sky130_fd_sc_hd__o21a_1 _10676_ (.A1(\sa_inst.cols_l2a:1.l2a_i._09_[6] ),
    .A2(_04591_),
    .B1(_04594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00010_));
 sky130_fd_sc_hd__buf_2 _10677_ (.A(\sa_inst.sak._10_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04595_));
 sky130_fd_sc_hd__clkbuf_1 _10678_ (.A(_04595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04596_));
 sky130_fd_sc_hd__and2_1 _10679_ (.A(_01057_),
    .B(_04596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04597_));
 sky130_fd_sc_hd__clkbuf_1 _10680_ (.A(_04597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00011_));
 sky130_fd_sc_hd__and2_1 _10681_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[1] ),
    .B(_04596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04598_));
 sky130_fd_sc_hd__clkbuf_1 _10682_ (.A(_04598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00012_));
 sky130_fd_sc_hd__and2_1 _10683_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[2] ),
    .B(_04596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04599_));
 sky130_fd_sc_hd__clkbuf_1 _10684_ (.A(_04599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00013_));
 sky130_fd_sc_hd__and2_1 _10685_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[3] ),
    .B(_04596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04600_));
 sky130_fd_sc_hd__clkbuf_1 _10686_ (.A(_04600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00014_));
 sky130_fd_sc_hd__and2_1 _10687_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[4] ),
    .B(_04596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04601_));
 sky130_fd_sc_hd__clkbuf_1 _10688_ (.A(_04601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00015_));
 sky130_fd_sc_hd__clkbuf_1 _10689_ (.A(_04595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04602_));
 sky130_fd_sc_hd__and2_1 _10690_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[5] ),
    .B(_04602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04603_));
 sky130_fd_sc_hd__clkbuf_1 _10691_ (.A(_04603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00016_));
 sky130_fd_sc_hd__and2_1 _10692_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[6] ),
    .B(_04602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04604_));
 sky130_fd_sc_hd__clkbuf_1 _10693_ (.A(_04604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00017_));
 sky130_fd_sc_hd__and2_1 _10694_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[7] ),
    .B(_04602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04605_));
 sky130_fd_sc_hd__clkbuf_1 _10695_ (.A(_04605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00018_));
 sky130_fd_sc_hd__and2_1 _10696_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[8] ),
    .B(_04602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04606_));
 sky130_fd_sc_hd__clkbuf_1 _10697_ (.A(_04606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00019_));
 sky130_fd_sc_hd__and2_1 _10698_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[9] ),
    .B(_04602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04607_));
 sky130_fd_sc_hd__clkbuf_1 _10699_ (.A(_04607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00020_));
 sky130_fd_sc_hd__clkbuf_1 _10700_ (.A(\sa_inst.sak._10_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04608_));
 sky130_fd_sc_hd__and2_1 _10701_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[10] ),
    .B(_04608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04609_));
 sky130_fd_sc_hd__clkbuf_1 _10702_ (.A(_04609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00021_));
 sky130_fd_sc_hd__and2_1 _10703_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[11] ),
    .B(_04608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04610_));
 sky130_fd_sc_hd__clkbuf_1 _10704_ (.A(_04610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00022_));
 sky130_fd_sc_hd__and2_1 _10705_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[12] ),
    .B(_04608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04611_));
 sky130_fd_sc_hd__clkbuf_1 _10706_ (.A(_04611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00023_));
 sky130_fd_sc_hd__and2_1 _10707_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[13] ),
    .B(_04608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04612_));
 sky130_fd_sc_hd__clkbuf_1 _10708_ (.A(_04612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00024_));
 sky130_fd_sc_hd__and2_1 _10709_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[14] ),
    .B(_04608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04613_));
 sky130_fd_sc_hd__clkbuf_1 _10710_ (.A(_04613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00025_));
 sky130_fd_sc_hd__clkbuf_1 _10711_ (.A(\sa_inst.sak._10_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04614_));
 sky130_fd_sc_hd__and2_1 _10712_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[15] ),
    .B(_04614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04615_));
 sky130_fd_sc_hd__clkbuf_1 _10713_ (.A(_04615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00026_));
 sky130_fd_sc_hd__and2_1 _10714_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[16] ),
    .B(_04614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04616_));
 sky130_fd_sc_hd__clkbuf_1 _10715_ (.A(_04616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00027_));
 sky130_fd_sc_hd__and2_1 _10716_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[17] ),
    .B(_04614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04617_));
 sky130_fd_sc_hd__clkbuf_1 _10717_ (.A(_04617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00028_));
 sky130_fd_sc_hd__and2_1 _10718_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[18] ),
    .B(_04614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04618_));
 sky130_fd_sc_hd__clkbuf_1 _10719_ (.A(_04618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00029_));
 sky130_fd_sc_hd__and2_1 _10720_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[19] ),
    .B(_04614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04619_));
 sky130_fd_sc_hd__clkbuf_1 _10721_ (.A(_04619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00030_));
 sky130_fd_sc_hd__clkbuf_1 _10722_ (.A(\sa_inst.sak._10_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04620_));
 sky130_fd_sc_hd__and2_1 _10723_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[20] ),
    .B(_04620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04621_));
 sky130_fd_sc_hd__clkbuf_1 _10724_ (.A(_04621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00031_));
 sky130_fd_sc_hd__and2_1 _10725_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[21] ),
    .B(_04620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04622_));
 sky130_fd_sc_hd__clkbuf_1 _10726_ (.A(_04622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00032_));
 sky130_fd_sc_hd__and2_1 _10727_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[22] ),
    .B(_04620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04623_));
 sky130_fd_sc_hd__clkbuf_1 _10728_ (.A(_04623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00033_));
 sky130_fd_sc_hd__and2_1 _10729_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[23] ),
    .B(_04620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04624_));
 sky130_fd_sc_hd__clkbuf_1 _10730_ (.A(_04624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00034_));
 sky130_fd_sc_hd__and2_1 _10731_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[24] ),
    .B(_04620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04625_));
 sky130_fd_sc_hd__clkbuf_1 _10732_ (.A(_04625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00035_));
 sky130_fd_sc_hd__clkbuf_1 _10733_ (.A(\sa_inst.sak._10_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04626_));
 sky130_fd_sc_hd__and2_1 _10734_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[25] ),
    .B(_04626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04627_));
 sky130_fd_sc_hd__clkbuf_1 _10735_ (.A(_04627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00036_));
 sky130_fd_sc_hd__and2_1 _10736_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[26] ),
    .B(_04626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04628_));
 sky130_fd_sc_hd__clkbuf_1 _10737_ (.A(_04628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00037_));
 sky130_fd_sc_hd__and2_1 _10738_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[27] ),
    .B(_04626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04629_));
 sky130_fd_sc_hd__clkbuf_1 _10739_ (.A(_04629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00038_));
 sky130_fd_sc_hd__and2_1 _10740_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[28] ),
    .B(_04626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04630_));
 sky130_fd_sc_hd__clkbuf_1 _10741_ (.A(_04630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00039_));
 sky130_fd_sc_hd__and2_1 _10742_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[29] ),
    .B(_04626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04631_));
 sky130_fd_sc_hd__clkbuf_1 _10743_ (.A(_04631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00040_));
 sky130_fd_sc_hd__and2_1 _10744_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[30] ),
    .B(_04595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04632_));
 sky130_fd_sc_hd__clkbuf_1 _10745_ (.A(_04632_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00041_));
 sky130_fd_sc_hd__and2_1 _10746_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[31] ),
    .B(_04595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04633_));
 sky130_fd_sc_hd__clkbuf_1 _10747_ (.A(_04633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00042_));
 sky130_fd_sc_hd__and2_1 _10748_ (.A(\sa_inst.sak.rows:1.cols:1.pe_ij._02_ ),
    .B(_04595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04634_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10749_ (.A(_04634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00043_));
 sky130_fd_sc_hd__clkbuf_2 _10750_ (.A(_02580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04635_));
 sky130_fd_sc_hd__and2_1 _10751_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[0] ),
    .B(_04635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04636_));
 sky130_fd_sc_hd__clkbuf_1 _10752_ (.A(_04636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00044_));
 sky130_fd_sc_hd__and2_1 _10753_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[1] ),
    .B(_04635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04637_));
 sky130_fd_sc_hd__clkbuf_1 _10754_ (.A(_04637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00045_));
 sky130_fd_sc_hd__and2_1 _10755_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[2] ),
    .B(_04635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04638_));
 sky130_fd_sc_hd__clkbuf_1 _10756_ (.A(_04638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00046_));
 sky130_fd_sc_hd__and2_1 _10757_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[3] ),
    .B(_04635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04639_));
 sky130_fd_sc_hd__clkbuf_1 _10758_ (.A(_04639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00047_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10759_ (.A(_02580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04640_));
 sky130_fd_sc_hd__and2_1 _10760_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[4] ),
    .B(_04640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04641_));
 sky130_fd_sc_hd__clkbuf_1 _10761_ (.A(_04641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00048_));
 sky130_fd_sc_hd__and2_1 _10762_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[5] ),
    .B(_04640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04642_));
 sky130_fd_sc_hd__clkbuf_1 _10763_ (.A(_04642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00049_));
 sky130_fd_sc_hd__and2_1 _10764_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[6] ),
    .B(_04640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04643_));
 sky130_fd_sc_hd__clkbuf_1 _10765_ (.A(_04643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00050_));
 sky130_fd_sc_hd__and2_1 _10766_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[7] ),
    .B(_04640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04644_));
 sky130_fd_sc_hd__clkbuf_1 _10767_ (.A(_04644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00051_));
 sky130_fd_sc_hd__and2_1 _10768_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[8] ),
    .B(_04640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04645_));
 sky130_fd_sc_hd__clkbuf_1 _10769_ (.A(_04645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00052_));
 sky130_fd_sc_hd__clkbuf_1 _10770_ (.A(_02580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04646_));
 sky130_fd_sc_hd__and2_1 _10771_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[9] ),
    .B(_04646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04647_));
 sky130_fd_sc_hd__clkbuf_1 _10772_ (.A(_04647_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00053_));
 sky130_fd_sc_hd__and2_1 _10773_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[10] ),
    .B(_04646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04648_));
 sky130_fd_sc_hd__clkbuf_1 _10774_ (.A(_04648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00054_));
 sky130_fd_sc_hd__and2_1 _10775_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[11] ),
    .B(_04646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04649_));
 sky130_fd_sc_hd__clkbuf_1 _10776_ (.A(_04649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00055_));
 sky130_fd_sc_hd__and2_1 _10777_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[12] ),
    .B(_04646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04650_));
 sky130_fd_sc_hd__clkbuf_1 _10778_ (.A(_04650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00056_));
 sky130_fd_sc_hd__and2_1 _10779_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[13] ),
    .B(_04646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04651_));
 sky130_fd_sc_hd__clkbuf_1 _10780_ (.A(_04651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00057_));
 sky130_fd_sc_hd__clkbuf_1 _10781_ (.A(_02580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04652_));
 sky130_fd_sc_hd__and2_1 _10782_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[14] ),
    .B(_04652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04653_));
 sky130_fd_sc_hd__clkbuf_1 _10783_ (.A(_04653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00058_));
 sky130_fd_sc_hd__and2_1 _10784_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[15] ),
    .B(_04652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04654_));
 sky130_fd_sc_hd__clkbuf_1 _10785_ (.A(_04654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00059_));
 sky130_fd_sc_hd__and2_1 _10786_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[16] ),
    .B(_04652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04655_));
 sky130_fd_sc_hd__clkbuf_1 _10787_ (.A(_04655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00060_));
 sky130_fd_sc_hd__and2_1 _10788_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[17] ),
    .B(_04652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04656_));
 sky130_fd_sc_hd__clkbuf_1 _10789_ (.A(_04656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00061_));
 sky130_fd_sc_hd__and2_1 _10790_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[18] ),
    .B(_04652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04657_));
 sky130_fd_sc_hd__clkbuf_1 _10791_ (.A(_04657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00062_));
 sky130_fd_sc_hd__clkbuf_1 _10792_ (.A(_02543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04658_));
 sky130_fd_sc_hd__and2_1 _10793_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[19] ),
    .B(_04658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04659_));
 sky130_fd_sc_hd__clkbuf_1 _10794_ (.A(_04659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00063_));
 sky130_fd_sc_hd__and2_1 _10795_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[20] ),
    .B(_04658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04660_));
 sky130_fd_sc_hd__clkbuf_1 _10796_ (.A(_04660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00064_));
 sky130_fd_sc_hd__and2_1 _10797_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[21] ),
    .B(_04658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04661_));
 sky130_fd_sc_hd__clkbuf_1 _10798_ (.A(_04661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00065_));
 sky130_fd_sc_hd__and2_1 _10799_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[22] ),
    .B(_04658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04662_));
 sky130_fd_sc_hd__clkbuf_1 _10800_ (.A(_04662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00066_));
 sky130_fd_sc_hd__and2_1 _10801_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[23] ),
    .B(_04658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04663_));
 sky130_fd_sc_hd__clkbuf_1 _10802_ (.A(_04663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00067_));
 sky130_fd_sc_hd__clkbuf_1 _10803_ (.A(_02543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04664_));
 sky130_fd_sc_hd__and2_1 _10804_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[24] ),
    .B(_04664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04665_));
 sky130_fd_sc_hd__clkbuf_1 _10805_ (.A(_04665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00068_));
 sky130_fd_sc_hd__and2_1 _10806_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[25] ),
    .B(_04664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04666_));
 sky130_fd_sc_hd__clkbuf_1 _10807_ (.A(_04666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00069_));
 sky130_fd_sc_hd__and2_1 _10808_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[26] ),
    .B(_04664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04667_));
 sky130_fd_sc_hd__clkbuf_1 _10809_ (.A(_04667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00070_));
 sky130_fd_sc_hd__and2_1 _10810_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[27] ),
    .B(_04664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04668_));
 sky130_fd_sc_hd__clkbuf_1 _10811_ (.A(_04668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00071_));
 sky130_fd_sc_hd__and2_1 _10812_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[28] ),
    .B(_04664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04669_));
 sky130_fd_sc_hd__clkbuf_1 _10813_ (.A(_04669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00072_));
 sky130_fd_sc_hd__and2_1 _10814_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[29] ),
    .B(_02540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04670_));
 sky130_fd_sc_hd__clkbuf_1 _10815_ (.A(_04670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00073_));
 sky130_fd_sc_hd__and2_1 _10816_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[30] ),
    .B(_02540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04671_));
 sky130_fd_sc_hd__clkbuf_1 _10817_ (.A(_04671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00074_));
 sky130_fd_sc_hd__and2_1 _10818_ (.A(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[31] ),
    .B(_02540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04672_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10819_ (.A(_04672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00075_));
 sky130_fd_sc_hd__and2_1 _10820_ (.A(_04635_),
    .B(\sa_inst.sak.rows:1.cols:2.pe_ij._02_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04673_));
 sky130_fd_sc_hd__clkbuf_1 _10821_ (.A(_04673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00076_));
 sky130_fd_sc_hd__buf_2 _10822_ (.A(_03634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04674_));
 sky130_fd_sc_hd__and2_1 _10823_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[0] ),
    .B(_04674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04675_));
 sky130_fd_sc_hd__clkbuf_1 _10824_ (.A(_04675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00077_));
 sky130_fd_sc_hd__and2_1 _10825_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[1] ),
    .B(_04674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04676_));
 sky130_fd_sc_hd__clkbuf_1 _10826_ (.A(_04676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00078_));
 sky130_fd_sc_hd__and2_1 _10827_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[2] ),
    .B(_04674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04677_));
 sky130_fd_sc_hd__clkbuf_1 _10828_ (.A(_04677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00079_));
 sky130_fd_sc_hd__and2_1 _10829_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[3] ),
    .B(_04674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04678_));
 sky130_fd_sc_hd__clkbuf_1 _10830_ (.A(_04678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00080_));
 sky130_fd_sc_hd__clkbuf_2 _10831_ (.A(_02796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04679_));
 sky130_fd_sc_hd__clkbuf_1 _10832_ (.A(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04680_));
 sky130_fd_sc_hd__and2_1 _10833_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[4] ),
    .B(_04680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04681_));
 sky130_fd_sc_hd__clkbuf_1 _10834_ (.A(_04681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00081_));
 sky130_fd_sc_hd__and2_1 _10835_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[5] ),
    .B(_04680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04682_));
 sky130_fd_sc_hd__clkbuf_1 _10836_ (.A(_04682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00082_));
 sky130_fd_sc_hd__and2_1 _10837_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[6] ),
    .B(_04680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04683_));
 sky130_fd_sc_hd__clkbuf_1 _10838_ (.A(_04683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00083_));
 sky130_fd_sc_hd__and2_1 _10839_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[7] ),
    .B(_04680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04684_));
 sky130_fd_sc_hd__clkbuf_1 _10840_ (.A(_04684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00084_));
 sky130_fd_sc_hd__and2_1 _10841_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[8] ),
    .B(_04680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04685_));
 sky130_fd_sc_hd__clkbuf_1 _10842_ (.A(_04685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00085_));
 sky130_fd_sc_hd__clkbuf_1 _10843_ (.A(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04686_));
 sky130_fd_sc_hd__and2_1 _10844_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[9] ),
    .B(_04686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04687_));
 sky130_fd_sc_hd__clkbuf_1 _10845_ (.A(_04687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00086_));
 sky130_fd_sc_hd__and2_1 _10846_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[10] ),
    .B(_04686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04688_));
 sky130_fd_sc_hd__clkbuf_1 _10847_ (.A(_04688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00087_));
 sky130_fd_sc_hd__and2_1 _10848_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[11] ),
    .B(_04686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04689_));
 sky130_fd_sc_hd__clkbuf_1 _10849_ (.A(_04689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00088_));
 sky130_fd_sc_hd__and2_1 _10850_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[12] ),
    .B(_04686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04690_));
 sky130_fd_sc_hd__clkbuf_1 _10851_ (.A(_04690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00089_));
 sky130_fd_sc_hd__and2_1 _10852_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[13] ),
    .B(_04686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04691_));
 sky130_fd_sc_hd__clkbuf_1 _10853_ (.A(_04691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00090_));
 sky130_fd_sc_hd__clkbuf_1 _10854_ (.A(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04692_));
 sky130_fd_sc_hd__and2_1 _10855_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[14] ),
    .B(_04692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04693_));
 sky130_fd_sc_hd__clkbuf_1 _10856_ (.A(_04693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00091_));
 sky130_fd_sc_hd__and2_1 _10857_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[15] ),
    .B(_04692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04694_));
 sky130_fd_sc_hd__clkbuf_1 _10858_ (.A(_04694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00092_));
 sky130_fd_sc_hd__and2_1 _10859_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[16] ),
    .B(_04692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04695_));
 sky130_fd_sc_hd__clkbuf_1 _10860_ (.A(_04695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00093_));
 sky130_fd_sc_hd__and2_1 _10861_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[17] ),
    .B(_04692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04696_));
 sky130_fd_sc_hd__clkbuf_1 _10862_ (.A(_04696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00094_));
 sky130_fd_sc_hd__and2_1 _10863_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[18] ),
    .B(_04692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04697_));
 sky130_fd_sc_hd__clkbuf_1 _10864_ (.A(_04697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00095_));
 sky130_fd_sc_hd__clkbuf_1 _10865_ (.A(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04698_));
 sky130_fd_sc_hd__and2_1 _10866_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[19] ),
    .B(_04698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04699_));
 sky130_fd_sc_hd__clkbuf_1 _10867_ (.A(_04699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00096_));
 sky130_fd_sc_hd__and2_1 _10868_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[20] ),
    .B(_04698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04700_));
 sky130_fd_sc_hd__clkbuf_1 _10869_ (.A(_04700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00097_));
 sky130_fd_sc_hd__and2_1 _10870_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[21] ),
    .B(_04698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04701_));
 sky130_fd_sc_hd__clkbuf_1 _10871_ (.A(_04701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00098_));
 sky130_fd_sc_hd__and2_1 _10872_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[22] ),
    .B(_04698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04702_));
 sky130_fd_sc_hd__clkbuf_1 _10873_ (.A(_04702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00099_));
 sky130_fd_sc_hd__and2_1 _10874_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[23] ),
    .B(_04698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04703_));
 sky130_fd_sc_hd__clkbuf_1 _10875_ (.A(_04703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00100_));
 sky130_fd_sc_hd__clkbuf_1 _10876_ (.A(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04704_));
 sky130_fd_sc_hd__and2_1 _10877_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[24] ),
    .B(_04704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04705_));
 sky130_fd_sc_hd__clkbuf_1 _10878_ (.A(_04705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00101_));
 sky130_fd_sc_hd__and2_1 _10879_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[25] ),
    .B(_04704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04706_));
 sky130_fd_sc_hd__clkbuf_1 _10880_ (.A(_04706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00102_));
 sky130_fd_sc_hd__and2_1 _10881_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[26] ),
    .B(_04704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04707_));
 sky130_fd_sc_hd__clkbuf_1 _10882_ (.A(_04707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00103_));
 sky130_fd_sc_hd__and2_1 _10883_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[27] ),
    .B(_04704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04708_));
 sky130_fd_sc_hd__clkbuf_1 _10884_ (.A(_04708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00104_));
 sky130_fd_sc_hd__and2_1 _10885_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[28] ),
    .B(_04704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04709_));
 sky130_fd_sc_hd__clkbuf_1 _10886_ (.A(_04709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00105_));
 sky130_fd_sc_hd__and2_1 _10887_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[29] ),
    .B(_02797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04710_));
 sky130_fd_sc_hd__clkbuf_1 _10888_ (.A(_04710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00106_));
 sky130_fd_sc_hd__and2_1 _10889_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[30] ),
    .B(_02797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04711_));
 sky130_fd_sc_hd__clkbuf_1 _10890_ (.A(_04711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00107_));
 sky130_fd_sc_hd__and2_1 _10891_ (.A(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[31] ),
    .B(_02797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04712_));
 sky130_fd_sc_hd__clkbuf_1 _10892_ (.A(_04712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00108_));
 sky130_fd_sc_hd__and2_1 _10893_ (.A(_04674_),
    .B(\sa_inst.sak.rows:1.cols:3.pe_ij._02_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04713_));
 sky130_fd_sc_hd__clkbuf_1 _10894_ (.A(_04713_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00109_));
 sky130_fd_sc_hd__xor2_1 _10895_ (.A(\fifo_inst.mem.RD1_ADDR[3] ),
    .B(\fifo_inst.mem.WR1_ADDR[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04714_));
 sky130_fd_sc_hd__xor2_1 _10896_ (.A(\fifo_inst.mem.RD1_ADDR[0] ),
    .B(\fifo_inst.mem.WR1_ADDR[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04715_));
 sky130_fd_sc_hd__xor2_1 _10897_ (.A(\fifo_inst.mem.RD1_ADDR[1] ),
    .B(\fifo_inst.mem.WR1_ADDR[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04716_));
 sky130_fd_sc_hd__xor2_1 _10898_ (.A(\fifo_inst.mem.RD1_ADDR[2] ),
    .B(\fifo_inst.mem.WR1_ADDR[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04717_));
 sky130_fd_sc_hd__or4_1 _10899_ (.A(_04714_),
    .B(_04715_),
    .C(_04716_),
    .D(_04717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04718_));
 sky130_fd_sc_hd__xnor2_1 _10900_ (.A(\fifo_inst.rRdPtr[4] ),
    .B(\fifo_inst.rWrPtr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04719_));
 sky130_fd_sc_hd__or2b_1 _10901_ (.A(_04718_),
    .B_N(_04719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04720_));
 sky130_fd_sc_hd__inv_2 _10902_ (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04721_));
 sky130_fd_sc_hd__o21ai_1 _10903_ (.A1(_04721_),
    .A2(\fifo_inst.rEmpty ),
    .B1(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04722_));
 sky130_fd_sc_hd__o21a_1 _10904_ (.A1(net55),
    .A2(_04720_),
    .B1(_04722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04723_));
 sky130_fd_sc_hd__buf_2 _10905_ (.A(_04723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04724_));
 sky130_fd_sc_hd__buf_2 _10906_ (.A(_04724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04725_));
 sky130_fd_sc_hd__clkbuf_2 _10907_ (.A(_04725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04726_));
 sky130_fd_sc_hd__clkbuf_2 _10908_ (.A(\fifo_inst.mem.RD1_ADDR[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04727_));
 sky130_fd_sc_hd__buf_2 _10909_ (.A(_04727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04728_));
 sky130_fd_sc_hd__clkbuf_2 _10910_ (.A(_04728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04729_));
 sky130_fd_sc_hd__clkbuf_4 _10911_ (.A(\fifo_inst.mem.RD1_ADDR[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04730_));
 sky130_fd_sc_hd__clkbuf_4 _10912_ (.A(_04730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04731_));
 sky130_fd_sc_hd__buf_2 _10913_ (.A(_04731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04732_));
 sky130_fd_sc_hd__buf_2 _10914_ (.A(_04732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04733_));
 sky130_fd_sc_hd__clkbuf_2 _10915_ (.A(\fifo_inst.mem.RD1_ADDR[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04734_));
 sky130_fd_sc_hd__clkbuf_4 _10916_ (.A(_04734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04735_));
 sky130_fd_sc_hd__clkbuf_2 _10917_ (.A(_04735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04736_));
 sky130_fd_sc_hd__buf_2 _10918_ (.A(_04736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04737_));
 sky130_fd_sc_hd__mux4_1 _10919_ (.A0(\fifo_inst.mem.rMemory[8][0] ),
    .A1(\fifo_inst.mem.rMemory[9][0] ),
    .A2(\fifo_inst.mem.rMemory[10][0] ),
    .A3(\fifo_inst.mem.rMemory[11][0] ),
    .S0(_04733_),
    .S1(_04737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04738_));
 sky130_fd_sc_hd__buf_6 _10920_ (.A(\fifo_inst.mem.RD1_ADDR[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04739_));
 sky130_fd_sc_hd__buf_2 _10921_ (.A(_04739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04740_));
 sky130_fd_sc_hd__clkbuf_2 _10922_ (.A(_04735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04741_));
 sky130_fd_sc_hd__mux4_1 _10923_ (.A0(\fifo_inst.mem.rMemory[12][0] ),
    .A1(\fifo_inst.mem.rMemory[13][0] ),
    .A2(\fifo_inst.mem.rMemory[14][0] ),
    .A3(\fifo_inst.mem.rMemory[15][0] ),
    .S0(_04740_),
    .S1(_04741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04742_));
 sky130_fd_sc_hd__clkbuf_4 _10924_ (.A(_04727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04743_));
 sky130_fd_sc_hd__clkbuf_1 _10925_ (.A(_04743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04744_));
 sky130_fd_sc_hd__or2b_1 _10926_ (.A(_04742_),
    .B_N(_04744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04745_));
 sky130_fd_sc_hd__clkbuf_4 _10927_ (.A(\fifo_inst.mem.RD1_ADDR[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04746_));
 sky130_fd_sc_hd__clkbuf_2 _10928_ (.A(_04746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04747_));
 sky130_fd_sc_hd__clkbuf_2 _10929_ (.A(_04747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04748_));
 sky130_fd_sc_hd__o211a_1 _10930_ (.A1(_04729_),
    .A2(_04738_),
    .B1(_04745_),
    .C1(_04748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04749_));
 sky130_fd_sc_hd__clkbuf_4 _10931_ (.A(_04727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04750_));
 sky130_fd_sc_hd__clkbuf_2 _10932_ (.A(_04750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04751_));
 sky130_fd_sc_hd__buf_4 _10933_ (.A(\fifo_inst.mem.RD1_ADDR[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04752_));
 sky130_fd_sc_hd__buf_2 _10934_ (.A(_04752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04753_));
 sky130_fd_sc_hd__buf_4 _10935_ (.A(\fifo_inst.mem.RD1_ADDR[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04754_));
 sky130_fd_sc_hd__buf_2 _10936_ (.A(_04754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04755_));
 sky130_fd_sc_hd__mux4_1 _10937_ (.A0(\fifo_inst.mem.rMemory[4][0] ),
    .A1(\fifo_inst.mem.rMemory[5][0] ),
    .A2(\fifo_inst.mem.rMemory[6][0] ),
    .A3(\fifo_inst.mem.rMemory[7][0] ),
    .S0(_04753_),
    .S1(_04755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04756_));
 sky130_fd_sc_hd__inv_2 _10938_ (.A(_04756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04757_));
 sky130_fd_sc_hd__clkbuf_2 _10939_ (.A(_04743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04758_));
 sky130_fd_sc_hd__buf_2 _10940_ (.A(_04731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04759_));
 sky130_fd_sc_hd__buf_4 _10941_ (.A(_04734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04760_));
 sky130_fd_sc_hd__buf_2 _10942_ (.A(_04760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04761_));
 sky130_fd_sc_hd__mux4_1 _10943_ (.A0(\fifo_inst.mem.rMemory[0][0] ),
    .A1(\fifo_inst.mem.rMemory[1][0] ),
    .A2(\fifo_inst.mem.rMemory[2][0] ),
    .A3(\fifo_inst.mem.rMemory[3][0] ),
    .S0(_04759_),
    .S1(_04761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04762_));
 sky130_fd_sc_hd__nor2_1 _10944_ (.A(_04758_),
    .B(_04762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04763_));
 sky130_fd_sc_hd__buf_2 _10945_ (.A(_04746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04764_));
 sky130_fd_sc_hd__clkbuf_2 _10946_ (.A(_04764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04765_));
 sky130_fd_sc_hd__a211o_1 _10947_ (.A1(_04751_),
    .A2(_04757_),
    .B1(_04763_),
    .C1(_04765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04766_));
 sky130_fd_sc_hd__nand2_1 _10948_ (.A(_04766_),
    .B(_04725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04767_));
 sky130_fd_sc_hd__o22a_1 _10949_ (.A1(net30),
    .A2(_04726_),
    .B1(_04749_),
    .B2(_04767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00110_));
 sky130_fd_sc_hd__mux4_1 _10950_ (.A0(\fifo_inst.mem.rMemory[8][1] ),
    .A1(\fifo_inst.mem.rMemory[9][1] ),
    .A2(\fifo_inst.mem.rMemory[10][1] ),
    .A3(\fifo_inst.mem.rMemory[11][1] ),
    .S0(_04733_),
    .S1(_04737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04768_));
 sky130_fd_sc_hd__mux4_1 _10951_ (.A0(\fifo_inst.mem.rMemory[12][1] ),
    .A1(\fifo_inst.mem.rMemory[13][1] ),
    .A2(\fifo_inst.mem.rMemory[14][1] ),
    .A3(\fifo_inst.mem.rMemory[15][1] ),
    .S0(_04740_),
    .S1(_04741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04769_));
 sky130_fd_sc_hd__or2b_1 _10952_ (.A(_04769_),
    .B_N(_04744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04770_));
 sky130_fd_sc_hd__o211a_1 _10953_ (.A1(_04729_),
    .A2(_04768_),
    .B1(_04770_),
    .C1(_04748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04771_));
 sky130_fd_sc_hd__buf_2 _10954_ (.A(_04723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04772_));
 sky130_fd_sc_hd__buf_2 _10955_ (.A(_04772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04773_));
 sky130_fd_sc_hd__mux4_1 _10956_ (.A0(\fifo_inst.mem.rMemory[4][1] ),
    .A1(\fifo_inst.mem.rMemory[5][1] ),
    .A2(\fifo_inst.mem.rMemory[6][1] ),
    .A3(\fifo_inst.mem.rMemory[7][1] ),
    .S0(_04753_),
    .S1(_04755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04774_));
 sky130_fd_sc_hd__inv_2 _10957_ (.A(_04774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04775_));
 sky130_fd_sc_hd__clkbuf_2 _10958_ (.A(_04727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04776_));
 sky130_fd_sc_hd__mux4_1 _10959_ (.A0(\fifo_inst.mem.rMemory[0][1] ),
    .A1(\fifo_inst.mem.rMemory[1][1] ),
    .A2(\fifo_inst.mem.rMemory[2][1] ),
    .A3(\fifo_inst.mem.rMemory[3][1] ),
    .S0(_04759_),
    .S1(_04761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04777_));
 sky130_fd_sc_hd__nor2_1 _10960_ (.A(_04776_),
    .B(_04777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04778_));
 sky130_fd_sc_hd__a211o_1 _10961_ (.A1(_04751_),
    .A2(_04775_),
    .B1(_04778_),
    .C1(_04765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04779_));
 sky130_fd_sc_hd__nand2_1 _10962_ (.A(_04773_),
    .B(_04779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04780_));
 sky130_fd_sc_hd__o22a_1 _10963_ (.A1(net41),
    .A2(_04726_),
    .B1(_04771_),
    .B2(_04780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00111_));
 sky130_fd_sc_hd__mux4_1 _10964_ (.A0(\fifo_inst.mem.rMemory[8][2] ),
    .A1(\fifo_inst.mem.rMemory[9][2] ),
    .A2(\fifo_inst.mem.rMemory[10][2] ),
    .A3(\fifo_inst.mem.rMemory[11][2] ),
    .S0(_04733_),
    .S1(_04737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04781_));
 sky130_fd_sc_hd__mux4_1 _10965_ (.A0(\fifo_inst.mem.rMemory[12][2] ),
    .A1(\fifo_inst.mem.rMemory[13][2] ),
    .A2(\fifo_inst.mem.rMemory[14][2] ),
    .A3(\fifo_inst.mem.rMemory[15][2] ),
    .S0(_04740_),
    .S1(_04741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04782_));
 sky130_fd_sc_hd__or2b_1 _10966_ (.A(_04782_),
    .B_N(_04744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04783_));
 sky130_fd_sc_hd__o211a_1 _10967_ (.A1(_04729_),
    .A2(_04781_),
    .B1(_04783_),
    .C1(_04748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04784_));
 sky130_fd_sc_hd__buf_2 _10968_ (.A(_04772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04785_));
 sky130_fd_sc_hd__clkbuf_4 _10969_ (.A(_04730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04786_));
 sky130_fd_sc_hd__buf_2 _10970_ (.A(_04754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04787_));
 sky130_fd_sc_hd__mux4_1 _10971_ (.A0(\fifo_inst.mem.rMemory[4][2] ),
    .A1(\fifo_inst.mem.rMemory[5][2] ),
    .A2(\fifo_inst.mem.rMemory[6][2] ),
    .A3(\fifo_inst.mem.rMemory[7][2] ),
    .S0(_04786_),
    .S1(_04787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04788_));
 sky130_fd_sc_hd__inv_2 _10972_ (.A(_04788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04789_));
 sky130_fd_sc_hd__clkbuf_4 _10973_ (.A(\fifo_inst.mem.RD1_ADDR[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04790_));
 sky130_fd_sc_hd__buf_2 _10974_ (.A(_04790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04791_));
 sky130_fd_sc_hd__mux4_1 _10975_ (.A0(\fifo_inst.mem.rMemory[0][2] ),
    .A1(\fifo_inst.mem.rMemory[1][2] ),
    .A2(\fifo_inst.mem.rMemory[2][2] ),
    .A3(\fifo_inst.mem.rMemory[3][2] ),
    .S0(_04759_),
    .S1(_04761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04792_));
 sky130_fd_sc_hd__nor2_1 _10976_ (.A(_04791_),
    .B(_04792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04793_));
 sky130_fd_sc_hd__a211o_1 _10977_ (.A1(_04751_),
    .A2(_04789_),
    .B1(_04793_),
    .C1(_04765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04794_));
 sky130_fd_sc_hd__nand2_1 _10978_ (.A(_04785_),
    .B(_04794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04795_));
 sky130_fd_sc_hd__o22a_1 _10979_ (.A1(net46),
    .A2(_04726_),
    .B1(_04784_),
    .B2(_04795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00112_));
 sky130_fd_sc_hd__mux4_1 _10980_ (.A0(\fifo_inst.mem.rMemory[8][3] ),
    .A1(\fifo_inst.mem.rMemory[9][3] ),
    .A2(\fifo_inst.mem.rMemory[10][3] ),
    .A3(\fifo_inst.mem.rMemory[11][3] ),
    .S0(_04733_),
    .S1(_04737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04796_));
 sky130_fd_sc_hd__mux4_1 _10981_ (.A0(\fifo_inst.mem.rMemory[12][3] ),
    .A1(\fifo_inst.mem.rMemory[13][3] ),
    .A2(\fifo_inst.mem.rMemory[14][3] ),
    .A3(\fifo_inst.mem.rMemory[15][3] ),
    .S0(_04740_),
    .S1(_04741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04797_));
 sky130_fd_sc_hd__or2b_1 _10982_ (.A(_04797_),
    .B_N(_04744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04798_));
 sky130_fd_sc_hd__o211a_1 _10983_ (.A1(_04729_),
    .A2(_04796_),
    .B1(_04798_),
    .C1(_04748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04799_));
 sky130_fd_sc_hd__mux4_1 _10984_ (.A0(\fifo_inst.mem.rMemory[4][3] ),
    .A1(\fifo_inst.mem.rMemory[5][3] ),
    .A2(\fifo_inst.mem.rMemory[6][3] ),
    .A3(\fifo_inst.mem.rMemory[7][3] ),
    .S0(_04786_),
    .S1(_04787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04800_));
 sky130_fd_sc_hd__inv_2 _10985_ (.A(_04800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04801_));
 sky130_fd_sc_hd__mux4_1 _10986_ (.A0(\fifo_inst.mem.rMemory[0][3] ),
    .A1(\fifo_inst.mem.rMemory[1][3] ),
    .A2(\fifo_inst.mem.rMemory[2][3] ),
    .A3(\fifo_inst.mem.rMemory[3][3] ),
    .S0(_04759_),
    .S1(_04761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04802_));
 sky130_fd_sc_hd__nor2_1 _10987_ (.A(_04791_),
    .B(_04802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04803_));
 sky130_fd_sc_hd__a211o_1 _10988_ (.A1(_04751_),
    .A2(_04801_),
    .B1(_04803_),
    .C1(_04765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04804_));
 sky130_fd_sc_hd__nand2_1 _10989_ (.A(_04785_),
    .B(_04804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04805_));
 sky130_fd_sc_hd__o22a_1 _10990_ (.A1(net47),
    .A2(_04726_),
    .B1(_04799_),
    .B2(_04805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00113_));
 sky130_fd_sc_hd__buf_2 _10991_ (.A(_04728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04806_));
 sky130_fd_sc_hd__clkbuf_4 _10992_ (.A(_04739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04807_));
 sky130_fd_sc_hd__clkbuf_4 _10993_ (.A(_04807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04808_));
 sky130_fd_sc_hd__buf_2 _10994_ (.A(_04735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04809_));
 sky130_fd_sc_hd__buf_2 _10995_ (.A(_04809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04810_));
 sky130_fd_sc_hd__mux4_1 _10996_ (.A0(\fifo_inst.mem.rMemory[8][4] ),
    .A1(\fifo_inst.mem.rMemory[9][4] ),
    .A2(\fifo_inst.mem.rMemory[10][4] ),
    .A3(\fifo_inst.mem.rMemory[11][4] ),
    .S0(_04808_),
    .S1(_04810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04811_));
 sky130_fd_sc_hd__mux4_1 _10997_ (.A0(\fifo_inst.mem.rMemory[12][4] ),
    .A1(\fifo_inst.mem.rMemory[13][4] ),
    .A2(\fifo_inst.mem.rMemory[14][4] ),
    .A3(\fifo_inst.mem.rMemory[15][4] ),
    .S0(_04740_),
    .S1(_04741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04812_));
 sky130_fd_sc_hd__or2b_1 _10998_ (.A(_04812_),
    .B_N(_04744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04813_));
 sky130_fd_sc_hd__o211a_1 _10999_ (.A1(_04806_),
    .A2(_04811_),
    .B1(_04813_),
    .C1(_04748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04814_));
 sky130_fd_sc_hd__mux4_1 _11000_ (.A0(\fifo_inst.mem.rMemory[4][4] ),
    .A1(\fifo_inst.mem.rMemory[5][4] ),
    .A2(\fifo_inst.mem.rMemory[6][4] ),
    .A3(\fifo_inst.mem.rMemory[7][4] ),
    .S0(_04786_),
    .S1(_04787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04815_));
 sky130_fd_sc_hd__inv_2 _11001_ (.A(_04815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04816_));
 sky130_fd_sc_hd__mux4_1 _11002_ (.A0(\fifo_inst.mem.rMemory[0][4] ),
    .A1(\fifo_inst.mem.rMemory[1][4] ),
    .A2(\fifo_inst.mem.rMemory[2][4] ),
    .A3(\fifo_inst.mem.rMemory[3][4] ),
    .S0(_04759_),
    .S1(_04761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04817_));
 sky130_fd_sc_hd__nor2_1 _11003_ (.A(_04791_),
    .B(_04817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04818_));
 sky130_fd_sc_hd__a211o_1 _11004_ (.A1(_04751_),
    .A2(_04816_),
    .B1(_04818_),
    .C1(_04765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04819_));
 sky130_fd_sc_hd__nand2_1 _11005_ (.A(_04785_),
    .B(_04819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04820_));
 sky130_fd_sc_hd__o22a_1 _11006_ (.A1(net48),
    .A2(_04726_),
    .B1(_04814_),
    .B2(_04820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00114_));
 sky130_fd_sc_hd__clkbuf_4 _11007_ (.A(_04723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04821_));
 sky130_fd_sc_hd__clkbuf_2 _11008_ (.A(_04821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04822_));
 sky130_fd_sc_hd__mux4_1 _11009_ (.A0(\fifo_inst.mem.rMemory[8][5] ),
    .A1(\fifo_inst.mem.rMemory[9][5] ),
    .A2(\fifo_inst.mem.rMemory[10][5] ),
    .A3(\fifo_inst.mem.rMemory[11][5] ),
    .S0(_04808_),
    .S1(_04810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04823_));
 sky130_fd_sc_hd__buf_2 _11010_ (.A(_04752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04824_));
 sky130_fd_sc_hd__buf_2 _11011_ (.A(_04735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04825_));
 sky130_fd_sc_hd__mux4_1 _11012_ (.A0(\fifo_inst.mem.rMemory[12][5] ),
    .A1(\fifo_inst.mem.rMemory[13][5] ),
    .A2(\fifo_inst.mem.rMemory[14][5] ),
    .A3(\fifo_inst.mem.rMemory[15][5] ),
    .S0(_04824_),
    .S1(_04825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04826_));
 sky130_fd_sc_hd__clkbuf_1 _11013_ (.A(_04743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04827_));
 sky130_fd_sc_hd__or2b_1 _11014_ (.A(_04826_),
    .B_N(_04827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04828_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11015_ (.A(_04764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04829_));
 sky130_fd_sc_hd__o211a_1 _11016_ (.A1(_04806_),
    .A2(_04823_),
    .B1(_04828_),
    .C1(_04829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04830_));
 sky130_fd_sc_hd__clkbuf_2 _11017_ (.A(_04750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04831_));
 sky130_fd_sc_hd__mux4_1 _11018_ (.A0(\fifo_inst.mem.rMemory[4][5] ),
    .A1(\fifo_inst.mem.rMemory[5][5] ),
    .A2(\fifo_inst.mem.rMemory[6][5] ),
    .A3(\fifo_inst.mem.rMemory[7][5] ),
    .S0(_04786_),
    .S1(_04787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04832_));
 sky130_fd_sc_hd__inv_2 _11019_ (.A(_04832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04833_));
 sky130_fd_sc_hd__buf_2 _11020_ (.A(_04739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04834_));
 sky130_fd_sc_hd__clkbuf_2 _11021_ (.A(_04760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04835_));
 sky130_fd_sc_hd__mux4_1 _11022_ (.A0(\fifo_inst.mem.rMemory[0][5] ),
    .A1(\fifo_inst.mem.rMemory[1][5] ),
    .A2(\fifo_inst.mem.rMemory[2][5] ),
    .A3(\fifo_inst.mem.rMemory[3][5] ),
    .S0(_04834_),
    .S1(_04835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04836_));
 sky130_fd_sc_hd__nor2_1 _11023_ (.A(_04791_),
    .B(_04836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04837_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11024_ (.A(_04746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04838_));
 sky130_fd_sc_hd__a211o_1 _11025_ (.A1(_04831_),
    .A2(_04833_),
    .B1(_04837_),
    .C1(_04838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04839_));
 sky130_fd_sc_hd__nand2_1 _11026_ (.A(_04785_),
    .B(_04839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04840_));
 sky130_fd_sc_hd__o22a_1 _11027_ (.A1(net49),
    .A2(_04822_),
    .B1(_04830_),
    .B2(_04840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00115_));
 sky130_fd_sc_hd__mux4_1 _11028_ (.A0(\fifo_inst.mem.rMemory[8][6] ),
    .A1(\fifo_inst.mem.rMemory[9][6] ),
    .A2(\fifo_inst.mem.rMemory[10][6] ),
    .A3(\fifo_inst.mem.rMemory[11][6] ),
    .S0(_04808_),
    .S1(_04810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04841_));
 sky130_fd_sc_hd__mux4_1 _11029_ (.A0(\fifo_inst.mem.rMemory[12][6] ),
    .A1(\fifo_inst.mem.rMemory[13][6] ),
    .A2(\fifo_inst.mem.rMemory[14][6] ),
    .A3(\fifo_inst.mem.rMemory[15][6] ),
    .S0(_04824_),
    .S1(_04825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04842_));
 sky130_fd_sc_hd__or2b_1 _11030_ (.A(_04842_),
    .B_N(_04827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04843_));
 sky130_fd_sc_hd__o211a_1 _11031_ (.A1(_04806_),
    .A2(_04841_),
    .B1(_04843_),
    .C1(_04829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04844_));
 sky130_fd_sc_hd__mux4_1 _11032_ (.A0(\fifo_inst.mem.rMemory[4][6] ),
    .A1(\fifo_inst.mem.rMemory[5][6] ),
    .A2(\fifo_inst.mem.rMemory[6][6] ),
    .A3(\fifo_inst.mem.rMemory[7][6] ),
    .S0(_04786_),
    .S1(_04787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04845_));
 sky130_fd_sc_hd__inv_2 _11033_ (.A(_04845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04846_));
 sky130_fd_sc_hd__mux4_1 _11034_ (.A0(\fifo_inst.mem.rMemory[0][6] ),
    .A1(\fifo_inst.mem.rMemory[1][6] ),
    .A2(\fifo_inst.mem.rMemory[2][6] ),
    .A3(\fifo_inst.mem.rMemory[3][6] ),
    .S0(_04834_),
    .S1(_04835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04847_));
 sky130_fd_sc_hd__nor2_1 _11035_ (.A(_04791_),
    .B(_04847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04848_));
 sky130_fd_sc_hd__a211o_1 _11036_ (.A1(_04831_),
    .A2(_04846_),
    .B1(_04848_),
    .C1(_04838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04849_));
 sky130_fd_sc_hd__nand2_1 _11037_ (.A(_04785_),
    .B(_04849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04850_));
 sky130_fd_sc_hd__o22a_1 _11038_ (.A1(net50),
    .A2(_04822_),
    .B1(_04844_),
    .B2(_04850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00116_));
 sky130_fd_sc_hd__mux4_1 _11039_ (.A0(\fifo_inst.mem.rMemory[8][7] ),
    .A1(\fifo_inst.mem.rMemory[9][7] ),
    .A2(\fifo_inst.mem.rMemory[10][7] ),
    .A3(\fifo_inst.mem.rMemory[11][7] ),
    .S0(_04808_),
    .S1(_04810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04851_));
 sky130_fd_sc_hd__mux4_1 _11040_ (.A0(\fifo_inst.mem.rMemory[12][7] ),
    .A1(\fifo_inst.mem.rMemory[13][7] ),
    .A2(\fifo_inst.mem.rMemory[14][7] ),
    .A3(\fifo_inst.mem.rMemory[15][7] ),
    .S0(_04824_),
    .S1(_04825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04852_));
 sky130_fd_sc_hd__or2b_1 _11041_ (.A(_04852_),
    .B_N(_04827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04853_));
 sky130_fd_sc_hd__o211a_1 _11042_ (.A1(_04806_),
    .A2(_04851_),
    .B1(_04853_),
    .C1(_04829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04854_));
 sky130_fd_sc_hd__clkbuf_2 _11043_ (.A(_04772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04855_));
 sky130_fd_sc_hd__clkbuf_4 _11044_ (.A(_04730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04856_));
 sky130_fd_sc_hd__clkbuf_2 _11045_ (.A(_04754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04857_));
 sky130_fd_sc_hd__mux4_1 _11046_ (.A0(\fifo_inst.mem.rMemory[4][7] ),
    .A1(\fifo_inst.mem.rMemory[5][7] ),
    .A2(\fifo_inst.mem.rMemory[6][7] ),
    .A3(\fifo_inst.mem.rMemory[7][7] ),
    .S0(_04856_),
    .S1(_04857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04858_));
 sky130_fd_sc_hd__inv_2 _11047_ (.A(_04858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04859_));
 sky130_fd_sc_hd__clkbuf_2 _11048_ (.A(_04790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04860_));
 sky130_fd_sc_hd__mux4_1 _11049_ (.A0(\fifo_inst.mem.rMemory[0][7] ),
    .A1(\fifo_inst.mem.rMemory[1][7] ),
    .A2(\fifo_inst.mem.rMemory[2][7] ),
    .A3(\fifo_inst.mem.rMemory[3][7] ),
    .S0(_04834_),
    .S1(_04835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04861_));
 sky130_fd_sc_hd__nor2_1 _11050_ (.A(_04860_),
    .B(_04861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04862_));
 sky130_fd_sc_hd__a211o_1 _11051_ (.A1(_04831_),
    .A2(_04859_),
    .B1(_04862_),
    .C1(_04838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04863_));
 sky130_fd_sc_hd__nand2_1 _11052_ (.A(_04855_),
    .B(_04863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04864_));
 sky130_fd_sc_hd__o22a_1 _11053_ (.A1(net51),
    .A2(_04822_),
    .B1(_04854_),
    .B2(_04864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00117_));
 sky130_fd_sc_hd__mux4_1 _11054_ (.A0(\fifo_inst.mem.rMemory[8][8] ),
    .A1(\fifo_inst.mem.rMemory[9][8] ),
    .A2(\fifo_inst.mem.rMemory[10][8] ),
    .A3(\fifo_inst.mem.rMemory[11][8] ),
    .S0(_04808_),
    .S1(_04810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04865_));
 sky130_fd_sc_hd__mux4_1 _11055_ (.A0(\fifo_inst.mem.rMemory[12][8] ),
    .A1(\fifo_inst.mem.rMemory[13][8] ),
    .A2(\fifo_inst.mem.rMemory[14][8] ),
    .A3(\fifo_inst.mem.rMemory[15][8] ),
    .S0(_04824_),
    .S1(_04825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04866_));
 sky130_fd_sc_hd__or2b_1 _11056_ (.A(_04866_),
    .B_N(_04827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04867_));
 sky130_fd_sc_hd__o211a_1 _11057_ (.A1(_04806_),
    .A2(_04865_),
    .B1(_04867_),
    .C1(_04829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04868_));
 sky130_fd_sc_hd__mux4_1 _11058_ (.A0(\fifo_inst.mem.rMemory[4][8] ),
    .A1(\fifo_inst.mem.rMemory[5][8] ),
    .A2(\fifo_inst.mem.rMemory[6][8] ),
    .A3(\fifo_inst.mem.rMemory[7][8] ),
    .S0(_04856_),
    .S1(_04857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04869_));
 sky130_fd_sc_hd__inv_2 _11059_ (.A(_04869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04870_));
 sky130_fd_sc_hd__mux4_1 _11060_ (.A0(\fifo_inst.mem.rMemory[0][8] ),
    .A1(\fifo_inst.mem.rMemory[1][8] ),
    .A2(\fifo_inst.mem.rMemory[2][8] ),
    .A3(\fifo_inst.mem.rMemory[3][8] ),
    .S0(_04834_),
    .S1(_04835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04871_));
 sky130_fd_sc_hd__nor2_1 _11061_ (.A(_04860_),
    .B(_04871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04872_));
 sky130_fd_sc_hd__a211o_1 _11062_ (.A1(_04831_),
    .A2(_04870_),
    .B1(_04872_),
    .C1(_04838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04873_));
 sky130_fd_sc_hd__nand2_1 _11063_ (.A(_04855_),
    .B(_04873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04874_));
 sky130_fd_sc_hd__o22a_1 _11064_ (.A1(net52),
    .A2(_04822_),
    .B1(_04868_),
    .B2(_04874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00118_));
 sky130_fd_sc_hd__buf_2 _11065_ (.A(_04728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04875_));
 sky130_fd_sc_hd__clkbuf_4 _11066_ (.A(_04753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04876_));
 sky130_fd_sc_hd__buf_2 _11067_ (.A(_04755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04877_));
 sky130_fd_sc_hd__mux4_1 _11068_ (.A0(\fifo_inst.mem.rMemory[8][9] ),
    .A1(\fifo_inst.mem.rMemory[9][9] ),
    .A2(\fifo_inst.mem.rMemory[10][9] ),
    .A3(\fifo_inst.mem.rMemory[11][9] ),
    .S0(_04876_),
    .S1(_04877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04878_));
 sky130_fd_sc_hd__mux4_1 _11069_ (.A0(\fifo_inst.mem.rMemory[12][9] ),
    .A1(\fifo_inst.mem.rMemory[13][9] ),
    .A2(\fifo_inst.mem.rMemory[14][9] ),
    .A3(\fifo_inst.mem.rMemory[15][9] ),
    .S0(_04824_),
    .S1(_04825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04879_));
 sky130_fd_sc_hd__or2b_1 _11070_ (.A(_04879_),
    .B_N(_04827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04880_));
 sky130_fd_sc_hd__o211a_1 _11071_ (.A1(_04875_),
    .A2(_04878_),
    .B1(_04880_),
    .C1(_04829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04881_));
 sky130_fd_sc_hd__mux4_1 _11072_ (.A0(\fifo_inst.mem.rMemory[4][9] ),
    .A1(\fifo_inst.mem.rMemory[5][9] ),
    .A2(\fifo_inst.mem.rMemory[6][9] ),
    .A3(\fifo_inst.mem.rMemory[7][9] ),
    .S0(_04856_),
    .S1(_04857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04882_));
 sky130_fd_sc_hd__inv_2 _11073_ (.A(_04882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04883_));
 sky130_fd_sc_hd__mux4_1 _11074_ (.A0(\fifo_inst.mem.rMemory[0][9] ),
    .A1(\fifo_inst.mem.rMemory[1][9] ),
    .A2(\fifo_inst.mem.rMemory[2][9] ),
    .A3(\fifo_inst.mem.rMemory[3][9] ),
    .S0(_04834_),
    .S1(_04835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04884_));
 sky130_fd_sc_hd__nor2_1 _11075_ (.A(_04860_),
    .B(_04884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04885_));
 sky130_fd_sc_hd__a211o_1 _11076_ (.A1(_04831_),
    .A2(_04883_),
    .B1(_04885_),
    .C1(_04838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04886_));
 sky130_fd_sc_hd__nand2_1 _11077_ (.A(_04855_),
    .B(_04886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04887_));
 sky130_fd_sc_hd__o22a_1 _11078_ (.A1(net53),
    .A2(_04822_),
    .B1(_04881_),
    .B2(_04887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00119_));
 sky130_fd_sc_hd__buf_2 _11079_ (.A(_04821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04888_));
 sky130_fd_sc_hd__mux4_1 _11080_ (.A0(\fifo_inst.mem.rMemory[8][10] ),
    .A1(\fifo_inst.mem.rMemory[9][10] ),
    .A2(\fifo_inst.mem.rMemory[10][10] ),
    .A3(\fifo_inst.mem.rMemory[11][10] ),
    .S0(_04876_),
    .S1(_04877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04889_));
 sky130_fd_sc_hd__buf_2 _11081_ (.A(_04752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04890_));
 sky130_fd_sc_hd__clkbuf_2 _11082_ (.A(_04754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04891_));
 sky130_fd_sc_hd__mux4_1 _11083_ (.A0(\fifo_inst.mem.rMemory[12][10] ),
    .A1(\fifo_inst.mem.rMemory[13][10] ),
    .A2(\fifo_inst.mem.rMemory[14][10] ),
    .A3(\fifo_inst.mem.rMemory[15][10] ),
    .S0(_04890_),
    .S1(_04891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04892_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11084_ (.A(_04743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04893_));
 sky130_fd_sc_hd__or2b_1 _11085_ (.A(_04892_),
    .B_N(_04893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04894_));
 sky130_fd_sc_hd__clkbuf_2 _11086_ (.A(_04764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04895_));
 sky130_fd_sc_hd__o211a_1 _11087_ (.A1(_04875_),
    .A2(_04889_),
    .B1(_04894_),
    .C1(_04895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04896_));
 sky130_fd_sc_hd__clkbuf_2 _11088_ (.A(_04750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04897_));
 sky130_fd_sc_hd__mux4_1 _11089_ (.A0(\fifo_inst.mem.rMemory[4][10] ),
    .A1(\fifo_inst.mem.rMemory[5][10] ),
    .A2(\fifo_inst.mem.rMemory[6][10] ),
    .A3(\fifo_inst.mem.rMemory[7][10] ),
    .S0(_04856_),
    .S1(_04857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04898_));
 sky130_fd_sc_hd__inv_2 _11090_ (.A(_04898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04899_));
 sky130_fd_sc_hd__buf_2 _11091_ (.A(_04739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04900_));
 sky130_fd_sc_hd__clkbuf_2 _11092_ (.A(_04760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04901_));
 sky130_fd_sc_hd__mux4_1 _11093_ (.A0(\fifo_inst.mem.rMemory[0][10] ),
    .A1(\fifo_inst.mem.rMemory[1][10] ),
    .A2(\fifo_inst.mem.rMemory[2][10] ),
    .A3(\fifo_inst.mem.rMemory[3][10] ),
    .S0(_04900_),
    .S1(_04901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04902_));
 sky130_fd_sc_hd__nor2_1 _11094_ (.A(_04860_),
    .B(_04902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04903_));
 sky130_fd_sc_hd__clkbuf_2 _11095_ (.A(_04746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04904_));
 sky130_fd_sc_hd__a211o_1 _11096_ (.A1(_04897_),
    .A2(_04899_),
    .B1(_04903_),
    .C1(_04904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04905_));
 sky130_fd_sc_hd__nand2_1 _11097_ (.A(_04855_),
    .B(_04905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04906_));
 sky130_fd_sc_hd__o22a_1 _11098_ (.A1(net31),
    .A2(_04888_),
    .B1(_04896_),
    .B2(_04906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00120_));
 sky130_fd_sc_hd__mux4_1 _11099_ (.A0(\fifo_inst.mem.rMemory[8][11] ),
    .A1(\fifo_inst.mem.rMemory[9][11] ),
    .A2(\fifo_inst.mem.rMemory[10][11] ),
    .A3(\fifo_inst.mem.rMemory[11][11] ),
    .S0(_04876_),
    .S1(_04877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04907_));
 sky130_fd_sc_hd__mux4_1 _11100_ (.A0(\fifo_inst.mem.rMemory[12][11] ),
    .A1(\fifo_inst.mem.rMemory[13][11] ),
    .A2(\fifo_inst.mem.rMemory[14][11] ),
    .A3(\fifo_inst.mem.rMemory[15][11] ),
    .S0(_04890_),
    .S1(_04891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04908_));
 sky130_fd_sc_hd__or2b_1 _11101_ (.A(_04908_),
    .B_N(_04893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04909_));
 sky130_fd_sc_hd__o211a_1 _11102_ (.A1(_04875_),
    .A2(_04907_),
    .B1(_04909_),
    .C1(_04895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04910_));
 sky130_fd_sc_hd__mux4_1 _11103_ (.A0(\fifo_inst.mem.rMemory[4][11] ),
    .A1(\fifo_inst.mem.rMemory[5][11] ),
    .A2(\fifo_inst.mem.rMemory[6][11] ),
    .A3(\fifo_inst.mem.rMemory[7][11] ),
    .S0(_04856_),
    .S1(_04857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04911_));
 sky130_fd_sc_hd__inv_2 _11104_ (.A(_04911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04912_));
 sky130_fd_sc_hd__mux4_1 _11105_ (.A0(\fifo_inst.mem.rMemory[0][11] ),
    .A1(\fifo_inst.mem.rMemory[1][11] ),
    .A2(\fifo_inst.mem.rMemory[2][11] ),
    .A3(\fifo_inst.mem.rMemory[3][11] ),
    .S0(_04900_),
    .S1(_04901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04913_));
 sky130_fd_sc_hd__nor2_1 _11106_ (.A(_04860_),
    .B(_04913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04914_));
 sky130_fd_sc_hd__a211o_1 _11107_ (.A1(_04897_),
    .A2(_04912_),
    .B1(_04914_),
    .C1(_04904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04915_));
 sky130_fd_sc_hd__nand2_1 _11108_ (.A(_04855_),
    .B(_04915_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04916_));
 sky130_fd_sc_hd__o22a_1 _11109_ (.A1(net32),
    .A2(_04888_),
    .B1(_04910_),
    .B2(_04916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00121_));
 sky130_fd_sc_hd__mux4_1 _11110_ (.A0(\fifo_inst.mem.rMemory[8][12] ),
    .A1(\fifo_inst.mem.rMemory[9][12] ),
    .A2(\fifo_inst.mem.rMemory[10][12] ),
    .A3(\fifo_inst.mem.rMemory[11][12] ),
    .S0(_04876_),
    .S1(_04877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04917_));
 sky130_fd_sc_hd__mux4_1 _11111_ (.A0(\fifo_inst.mem.rMemory[12][12] ),
    .A1(\fifo_inst.mem.rMemory[13][12] ),
    .A2(\fifo_inst.mem.rMemory[14][12] ),
    .A3(\fifo_inst.mem.rMemory[15][12] ),
    .S0(_04890_),
    .S1(_04891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04918_));
 sky130_fd_sc_hd__or2b_1 _11112_ (.A(_04918_),
    .B_N(_04893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04919_));
 sky130_fd_sc_hd__o211a_1 _11113_ (.A1(_04875_),
    .A2(_04917_),
    .B1(_04919_),
    .C1(_04895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04920_));
 sky130_fd_sc_hd__clkbuf_4 _11114_ (.A(_04724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04921_));
 sky130_fd_sc_hd__buf_4 _11115_ (.A(_04730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04922_));
 sky130_fd_sc_hd__buf_4 _11116_ (.A(_04734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04923_));
 sky130_fd_sc_hd__mux4_1 _11117_ (.A0(\fifo_inst.mem.rMemory[4][12] ),
    .A1(\fifo_inst.mem.rMemory[5][12] ),
    .A2(\fifo_inst.mem.rMemory[6][12] ),
    .A3(\fifo_inst.mem.rMemory[7][12] ),
    .S0(_04922_),
    .S1(_04923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04924_));
 sky130_fd_sc_hd__inv_2 _11118_ (.A(_04924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04925_));
 sky130_fd_sc_hd__clkbuf_4 _11119_ (.A(_04790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04926_));
 sky130_fd_sc_hd__mux4_1 _11120_ (.A0(\fifo_inst.mem.rMemory[0][12] ),
    .A1(\fifo_inst.mem.rMemory[1][12] ),
    .A2(\fifo_inst.mem.rMemory[2][12] ),
    .A3(\fifo_inst.mem.rMemory[3][12] ),
    .S0(_04900_),
    .S1(_04901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04927_));
 sky130_fd_sc_hd__nor2_1 _11121_ (.A(_04926_),
    .B(_04927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04928_));
 sky130_fd_sc_hd__a211o_1 _11122_ (.A1(_04897_),
    .A2(_04925_),
    .B1(_04928_),
    .C1(_04904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04929_));
 sky130_fd_sc_hd__nand2_1 _11123_ (.A(_04921_),
    .B(_04929_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04930_));
 sky130_fd_sc_hd__o22a_1 _11124_ (.A1(net33),
    .A2(_04888_),
    .B1(_04920_),
    .B2(_04930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00122_));
 sky130_fd_sc_hd__mux4_1 _11125_ (.A0(\fifo_inst.mem.rMemory[8][13] ),
    .A1(\fifo_inst.mem.rMemory[9][13] ),
    .A2(\fifo_inst.mem.rMemory[10][13] ),
    .A3(\fifo_inst.mem.rMemory[11][13] ),
    .S0(_04876_),
    .S1(_04877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04931_));
 sky130_fd_sc_hd__mux4_1 _11126_ (.A0(\fifo_inst.mem.rMemory[12][13] ),
    .A1(\fifo_inst.mem.rMemory[13][13] ),
    .A2(\fifo_inst.mem.rMemory[14][13] ),
    .A3(\fifo_inst.mem.rMemory[15][13] ),
    .S0(_04890_),
    .S1(_04891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04932_));
 sky130_fd_sc_hd__or2b_1 _11127_ (.A(_04932_),
    .B_N(_04893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04933_));
 sky130_fd_sc_hd__o211a_1 _11128_ (.A1(_04875_),
    .A2(_04931_),
    .B1(_04933_),
    .C1(_04895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04934_));
 sky130_fd_sc_hd__mux4_1 _11129_ (.A0(\fifo_inst.mem.rMemory[4][13] ),
    .A1(\fifo_inst.mem.rMemory[5][13] ),
    .A2(\fifo_inst.mem.rMemory[6][13] ),
    .A3(\fifo_inst.mem.rMemory[7][13] ),
    .S0(_04922_),
    .S1(_04923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04935_));
 sky130_fd_sc_hd__inv_2 _11130_ (.A(_04935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04936_));
 sky130_fd_sc_hd__mux4_1 _11131_ (.A0(\fifo_inst.mem.rMemory[0][13] ),
    .A1(\fifo_inst.mem.rMemory[1][13] ),
    .A2(\fifo_inst.mem.rMemory[2][13] ),
    .A3(\fifo_inst.mem.rMemory[3][13] ),
    .S0(_04900_),
    .S1(_04901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04937_));
 sky130_fd_sc_hd__nor2_1 _11132_ (.A(_04926_),
    .B(_04937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04938_));
 sky130_fd_sc_hd__a211o_1 _11133_ (.A1(_04897_),
    .A2(_04936_),
    .B1(_04938_),
    .C1(_04904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04939_));
 sky130_fd_sc_hd__nand2_1 _11134_ (.A(_04921_),
    .B(_04939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04940_));
 sky130_fd_sc_hd__o22a_1 _11135_ (.A1(net34),
    .A2(_04888_),
    .B1(_04934_),
    .B2(_04940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00123_));
 sky130_fd_sc_hd__clkbuf_4 _11136_ (.A(_04750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04941_));
 sky130_fd_sc_hd__buf_4 _11137_ (.A(_04753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04942_));
 sky130_fd_sc_hd__buf_4 _11138_ (.A(_04755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04943_));
 sky130_fd_sc_hd__mux4_1 _11139_ (.A0(\fifo_inst.mem.rMemory[8][14] ),
    .A1(\fifo_inst.mem.rMemory[9][14] ),
    .A2(\fifo_inst.mem.rMemory[10][14] ),
    .A3(\fifo_inst.mem.rMemory[11][14] ),
    .S0(_04942_),
    .S1(_04943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04944_));
 sky130_fd_sc_hd__mux4_1 _11140_ (.A0(\fifo_inst.mem.rMemory[12][14] ),
    .A1(\fifo_inst.mem.rMemory[13][14] ),
    .A2(\fifo_inst.mem.rMemory[14][14] ),
    .A3(\fifo_inst.mem.rMemory[15][14] ),
    .S0(_04890_),
    .S1(_04891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04945_));
 sky130_fd_sc_hd__or2b_1 _11141_ (.A(_04945_),
    .B_N(_04893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04946_));
 sky130_fd_sc_hd__o211a_1 _11142_ (.A1(_04941_),
    .A2(_04944_),
    .B1(_04946_),
    .C1(_04895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04947_));
 sky130_fd_sc_hd__mux4_1 _11143_ (.A0(\fifo_inst.mem.rMemory[4][14] ),
    .A1(\fifo_inst.mem.rMemory[5][14] ),
    .A2(\fifo_inst.mem.rMemory[6][14] ),
    .A3(\fifo_inst.mem.rMemory[7][14] ),
    .S0(_04922_),
    .S1(_04923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04948_));
 sky130_fd_sc_hd__inv_2 _11144_ (.A(_04948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04949_));
 sky130_fd_sc_hd__mux4_1 _11145_ (.A0(\fifo_inst.mem.rMemory[0][14] ),
    .A1(\fifo_inst.mem.rMemory[1][14] ),
    .A2(\fifo_inst.mem.rMemory[2][14] ),
    .A3(\fifo_inst.mem.rMemory[3][14] ),
    .S0(_04900_),
    .S1(_04901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04950_));
 sky130_fd_sc_hd__nor2_1 _11146_ (.A(_04926_),
    .B(_04950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04951_));
 sky130_fd_sc_hd__a211o_1 _11147_ (.A1(_04897_),
    .A2(_04949_),
    .B1(_04951_),
    .C1(_04904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04952_));
 sky130_fd_sc_hd__nand2_1 _11148_ (.A(_04921_),
    .B(_04952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04953_));
 sky130_fd_sc_hd__o22a_1 _11149_ (.A1(net35),
    .A2(_04888_),
    .B1(_04947_),
    .B2(_04953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00124_));
 sky130_fd_sc_hd__clkbuf_2 _11150_ (.A(_04821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04954_));
 sky130_fd_sc_hd__mux4_1 _11151_ (.A0(\fifo_inst.mem.rMemory[8][15] ),
    .A1(\fifo_inst.mem.rMemory[9][15] ),
    .A2(\fifo_inst.mem.rMemory[10][15] ),
    .A3(\fifo_inst.mem.rMemory[11][15] ),
    .S0(_04942_),
    .S1(_04943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04955_));
 sky130_fd_sc_hd__clkbuf_4 _11152_ (.A(_04752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04956_));
 sky130_fd_sc_hd__buf_2 _11153_ (.A(_04754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04957_));
 sky130_fd_sc_hd__mux4_1 _11154_ (.A0(\fifo_inst.mem.rMemory[12][15] ),
    .A1(\fifo_inst.mem.rMemory[13][15] ),
    .A2(\fifo_inst.mem.rMemory[14][15] ),
    .A3(\fifo_inst.mem.rMemory[15][15] ),
    .S0(_04956_),
    .S1(_04957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04958_));
 sky130_fd_sc_hd__clkbuf_2 _11155_ (.A(_04743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04959_));
 sky130_fd_sc_hd__or2b_1 _11156_ (.A(_04958_),
    .B_N(_04959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04960_));
 sky130_fd_sc_hd__clkbuf_2 _11157_ (.A(_04764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04961_));
 sky130_fd_sc_hd__o211a_1 _11158_ (.A1(_04941_),
    .A2(_04955_),
    .B1(_04960_),
    .C1(_04961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04962_));
 sky130_fd_sc_hd__clkbuf_2 _11159_ (.A(_04790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04963_));
 sky130_fd_sc_hd__mux4_1 _11160_ (.A0(\fifo_inst.mem.rMemory[4][15] ),
    .A1(\fifo_inst.mem.rMemory[5][15] ),
    .A2(\fifo_inst.mem.rMemory[6][15] ),
    .A3(\fifo_inst.mem.rMemory[7][15] ),
    .S0(_04922_),
    .S1(_04923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04964_));
 sky130_fd_sc_hd__inv_2 _11161_ (.A(_04964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04965_));
 sky130_fd_sc_hd__buf_2 _11162_ (.A(_04739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04966_));
 sky130_fd_sc_hd__clkbuf_2 _11163_ (.A(_04735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04967_));
 sky130_fd_sc_hd__mux4_1 _11164_ (.A0(\fifo_inst.mem.rMemory[0][15] ),
    .A1(\fifo_inst.mem.rMemory[1][15] ),
    .A2(\fifo_inst.mem.rMemory[2][15] ),
    .A3(\fifo_inst.mem.rMemory[3][15] ),
    .S0(_04966_),
    .S1(_04967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04968_));
 sky130_fd_sc_hd__nor2_1 _11165_ (.A(_04926_),
    .B(_04968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04969_));
 sky130_fd_sc_hd__clkbuf_2 _11166_ (.A(_04746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04970_));
 sky130_fd_sc_hd__a211o_1 _11167_ (.A1(_04963_),
    .A2(_04965_),
    .B1(_04969_),
    .C1(_04970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04971_));
 sky130_fd_sc_hd__nand2_1 _11168_ (.A(_04921_),
    .B(_04971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04972_));
 sky130_fd_sc_hd__o22a_1 _11169_ (.A1(net36),
    .A2(_04954_),
    .B1(_04962_),
    .B2(_04972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00125_));
 sky130_fd_sc_hd__mux4_1 _11170_ (.A0(\fifo_inst.mem.rMemory[8][16] ),
    .A1(\fifo_inst.mem.rMemory[9][16] ),
    .A2(\fifo_inst.mem.rMemory[10][16] ),
    .A3(\fifo_inst.mem.rMemory[11][16] ),
    .S0(_04942_),
    .S1(_04943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04973_));
 sky130_fd_sc_hd__mux4_1 _11171_ (.A0(\fifo_inst.mem.rMemory[12][16] ),
    .A1(\fifo_inst.mem.rMemory[13][16] ),
    .A2(\fifo_inst.mem.rMemory[14][16] ),
    .A3(\fifo_inst.mem.rMemory[15][16] ),
    .S0(_04956_),
    .S1(_04957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04974_));
 sky130_fd_sc_hd__or2b_1 _11172_ (.A(_04974_),
    .B_N(_04959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04975_));
 sky130_fd_sc_hd__o211a_1 _11173_ (.A1(_04941_),
    .A2(_04973_),
    .B1(_04975_),
    .C1(_04961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04976_));
 sky130_fd_sc_hd__mux4_1 _11174_ (.A0(\fifo_inst.mem.rMemory[4][16] ),
    .A1(\fifo_inst.mem.rMemory[5][16] ),
    .A2(\fifo_inst.mem.rMemory[6][16] ),
    .A3(\fifo_inst.mem.rMemory[7][16] ),
    .S0(_04922_),
    .S1(_04923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04977_));
 sky130_fd_sc_hd__inv_2 _11175_ (.A(_04977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04978_));
 sky130_fd_sc_hd__mux4_1 _11176_ (.A0(\fifo_inst.mem.rMemory[0][16] ),
    .A1(\fifo_inst.mem.rMemory[1][16] ),
    .A2(\fifo_inst.mem.rMemory[2][16] ),
    .A3(\fifo_inst.mem.rMemory[3][16] ),
    .S0(_04966_),
    .S1(_04967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04979_));
 sky130_fd_sc_hd__nor2_1 _11177_ (.A(_04926_),
    .B(_04979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04980_));
 sky130_fd_sc_hd__a211o_1 _11178_ (.A1(_04963_),
    .A2(_04978_),
    .B1(_04980_),
    .C1(_04970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04981_));
 sky130_fd_sc_hd__nand2_1 _11179_ (.A(_04921_),
    .B(_04981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04982_));
 sky130_fd_sc_hd__o22a_1 _11180_ (.A1(net37),
    .A2(_04954_),
    .B1(_04976_),
    .B2(_04982_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00126_));
 sky130_fd_sc_hd__mux4_1 _11181_ (.A0(\fifo_inst.mem.rMemory[8][17] ),
    .A1(\fifo_inst.mem.rMemory[9][17] ),
    .A2(\fifo_inst.mem.rMemory[10][17] ),
    .A3(\fifo_inst.mem.rMemory[11][17] ),
    .S0(_04942_),
    .S1(_04943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04983_));
 sky130_fd_sc_hd__mux4_1 _11182_ (.A0(\fifo_inst.mem.rMemory[12][17] ),
    .A1(\fifo_inst.mem.rMemory[13][17] ),
    .A2(\fifo_inst.mem.rMemory[14][17] ),
    .A3(\fifo_inst.mem.rMemory[15][17] ),
    .S0(_04956_),
    .S1(_04957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04984_));
 sky130_fd_sc_hd__or2b_1 _11183_ (.A(_04984_),
    .B_N(_04959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04985_));
 sky130_fd_sc_hd__o211a_1 _11184_ (.A1(_04941_),
    .A2(_04983_),
    .B1(_04985_),
    .C1(_04961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04986_));
 sky130_fd_sc_hd__clkbuf_2 _11185_ (.A(_04724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04987_));
 sky130_fd_sc_hd__buf_2 _11186_ (.A(_04730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04988_));
 sky130_fd_sc_hd__clkbuf_2 _11187_ (.A(_04734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04989_));
 sky130_fd_sc_hd__mux4_1 _11188_ (.A0(\fifo_inst.mem.rMemory[4][17] ),
    .A1(\fifo_inst.mem.rMemory[5][17] ),
    .A2(\fifo_inst.mem.rMemory[6][17] ),
    .A3(\fifo_inst.mem.rMemory[7][17] ),
    .S0(_04988_),
    .S1(_04989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04990_));
 sky130_fd_sc_hd__inv_2 _11189_ (.A(_04990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04991_));
 sky130_fd_sc_hd__clkbuf_2 _11190_ (.A(_04790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04992_));
 sky130_fd_sc_hd__mux4_1 _11191_ (.A0(\fifo_inst.mem.rMemory[0][17] ),
    .A1(\fifo_inst.mem.rMemory[1][17] ),
    .A2(\fifo_inst.mem.rMemory[2][17] ),
    .A3(\fifo_inst.mem.rMemory[3][17] ),
    .S0(_04966_),
    .S1(_04967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04993_));
 sky130_fd_sc_hd__nor2_1 _11192_ (.A(_04992_),
    .B(_04993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04994_));
 sky130_fd_sc_hd__a211o_1 _11193_ (.A1(_04963_),
    .A2(_04991_),
    .B1(_04994_),
    .C1(_04970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04995_));
 sky130_fd_sc_hd__nand2_1 _11194_ (.A(_04987_),
    .B(_04995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04996_));
 sky130_fd_sc_hd__o22a_1 _11195_ (.A1(net38),
    .A2(_04954_),
    .B1(_04986_),
    .B2(_04996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00127_));
 sky130_fd_sc_hd__mux4_1 _11196_ (.A0(\fifo_inst.mem.rMemory[8][18] ),
    .A1(\fifo_inst.mem.rMemory[9][18] ),
    .A2(\fifo_inst.mem.rMemory[10][18] ),
    .A3(\fifo_inst.mem.rMemory[11][18] ),
    .S0(_04942_),
    .S1(_04943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04997_));
 sky130_fd_sc_hd__mux4_1 _11197_ (.A0(\fifo_inst.mem.rMemory[12][18] ),
    .A1(\fifo_inst.mem.rMemory[13][18] ),
    .A2(\fifo_inst.mem.rMemory[14][18] ),
    .A3(\fifo_inst.mem.rMemory[15][18] ),
    .S0(_04956_),
    .S1(_04957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04998_));
 sky130_fd_sc_hd__or2b_1 _11198_ (.A(_04998_),
    .B_N(_04959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04999_));
 sky130_fd_sc_hd__o211a_1 _11199_ (.A1(_04941_),
    .A2(_04997_),
    .B1(_04999_),
    .C1(_04961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05000_));
 sky130_fd_sc_hd__mux4_1 _11200_ (.A0(\fifo_inst.mem.rMemory[4][18] ),
    .A1(\fifo_inst.mem.rMemory[5][18] ),
    .A2(\fifo_inst.mem.rMemory[6][18] ),
    .A3(\fifo_inst.mem.rMemory[7][18] ),
    .S0(_04988_),
    .S1(_04989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05001_));
 sky130_fd_sc_hd__inv_2 _11201_ (.A(_05001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05002_));
 sky130_fd_sc_hd__mux4_1 _11202_ (.A0(\fifo_inst.mem.rMemory[0][18] ),
    .A1(\fifo_inst.mem.rMemory[1][18] ),
    .A2(\fifo_inst.mem.rMemory[2][18] ),
    .A3(\fifo_inst.mem.rMemory[3][18] ),
    .S0(_04966_),
    .S1(_04967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05003_));
 sky130_fd_sc_hd__nor2_1 _11203_ (.A(_04992_),
    .B(_05003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05004_));
 sky130_fd_sc_hd__a211o_1 _11204_ (.A1(_04963_),
    .A2(_05002_),
    .B1(_05004_),
    .C1(_04970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05005_));
 sky130_fd_sc_hd__nand2_1 _11205_ (.A(_04987_),
    .B(_05005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05006_));
 sky130_fd_sc_hd__o22a_1 _11206_ (.A1(net39),
    .A2(_04954_),
    .B1(_05000_),
    .B2(_05006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00128_));
 sky130_fd_sc_hd__clkbuf_4 _11207_ (.A(_04750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05007_));
 sky130_fd_sc_hd__clkbuf_4 _11208_ (.A(_04753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05008_));
 sky130_fd_sc_hd__buf_2 _11209_ (.A(_04755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05009_));
 sky130_fd_sc_hd__mux4_1 _11210_ (.A0(\fifo_inst.mem.rMemory[8][19] ),
    .A1(\fifo_inst.mem.rMemory[9][19] ),
    .A2(\fifo_inst.mem.rMemory[10][19] ),
    .A3(\fifo_inst.mem.rMemory[11][19] ),
    .S0(_05008_),
    .S1(_05009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05010_));
 sky130_fd_sc_hd__mux4_1 _11211_ (.A0(\fifo_inst.mem.rMemory[12][19] ),
    .A1(\fifo_inst.mem.rMemory[13][19] ),
    .A2(\fifo_inst.mem.rMemory[14][19] ),
    .A3(\fifo_inst.mem.rMemory[15][19] ),
    .S0(_04956_),
    .S1(_04957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05011_));
 sky130_fd_sc_hd__or2b_1 _11212_ (.A(_05011_),
    .B_N(_04959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05012_));
 sky130_fd_sc_hd__o211a_1 _11213_ (.A1(_05007_),
    .A2(_05010_),
    .B1(_05012_),
    .C1(_04961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05013_));
 sky130_fd_sc_hd__mux4_1 _11214_ (.A0(\fifo_inst.mem.rMemory[4][19] ),
    .A1(\fifo_inst.mem.rMemory[5][19] ),
    .A2(\fifo_inst.mem.rMemory[6][19] ),
    .A3(\fifo_inst.mem.rMemory[7][19] ),
    .S0(_04988_),
    .S1(_04989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05014_));
 sky130_fd_sc_hd__inv_2 _11215_ (.A(_05014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05015_));
 sky130_fd_sc_hd__mux4_1 _11216_ (.A0(\fifo_inst.mem.rMemory[0][19] ),
    .A1(\fifo_inst.mem.rMemory[1][19] ),
    .A2(\fifo_inst.mem.rMemory[2][19] ),
    .A3(\fifo_inst.mem.rMemory[3][19] ),
    .S0(_04966_),
    .S1(_04967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05016_));
 sky130_fd_sc_hd__nor2_1 _11217_ (.A(_04992_),
    .B(_05016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05017_));
 sky130_fd_sc_hd__a211o_1 _11218_ (.A1(_04963_),
    .A2(_05015_),
    .B1(_05017_),
    .C1(_04970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05018_));
 sky130_fd_sc_hd__nand2_1 _11219_ (.A(_04987_),
    .B(_05018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05019_));
 sky130_fd_sc_hd__o22a_1 _11220_ (.A1(net40),
    .A2(_04954_),
    .B1(_05013_),
    .B2(_05019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00129_));
 sky130_fd_sc_hd__mux4_1 _11221_ (.A0(\fifo_inst.mem.rMemory[8][20] ),
    .A1(\fifo_inst.mem.rMemory[9][20] ),
    .A2(\fifo_inst.mem.rMemory[10][20] ),
    .A3(\fifo_inst.mem.rMemory[11][20] ),
    .S0(_05008_),
    .S1(_05009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05020_));
 sky130_fd_sc_hd__mux4_1 _11222_ (.A0(\fifo_inst.mem.rMemory[12][20] ),
    .A1(\fifo_inst.mem.rMemory[13][20] ),
    .A2(\fifo_inst.mem.rMemory[14][20] ),
    .A3(\fifo_inst.mem.rMemory[15][20] ),
    .S0(_04807_),
    .S1(_04809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05021_));
 sky130_fd_sc_hd__or2b_1 _11223_ (.A(_05021_),
    .B_N(_04776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05022_));
 sky130_fd_sc_hd__buf_2 _11224_ (.A(_04764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05023_));
 sky130_fd_sc_hd__o211a_1 _11225_ (.A1(_05007_),
    .A2(_05020_),
    .B1(_05022_),
    .C1(_05023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05024_));
 sky130_fd_sc_hd__mux4_1 _11226_ (.A0(\fifo_inst.mem.rMemory[4][20] ),
    .A1(\fifo_inst.mem.rMemory[5][20] ),
    .A2(\fifo_inst.mem.rMemory[6][20] ),
    .A3(\fifo_inst.mem.rMemory[7][20] ),
    .S0(_04988_),
    .S1(_04989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05025_));
 sky130_fd_sc_hd__inv_2 _11227_ (.A(_05025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05026_));
 sky130_fd_sc_hd__mux4_1 _11228_ (.A0(\fifo_inst.mem.rMemory[0][20] ),
    .A1(\fifo_inst.mem.rMemory[1][20] ),
    .A2(\fifo_inst.mem.rMemory[2][20] ),
    .A3(\fifo_inst.mem.rMemory[3][20] ),
    .S0(_04732_),
    .S1(_04736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05027_));
 sky130_fd_sc_hd__nor2_1 _11229_ (.A(_04992_),
    .B(_05027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05028_));
 sky130_fd_sc_hd__a211o_1 _11230_ (.A1(_04758_),
    .A2(_05026_),
    .B1(_05028_),
    .C1(_04747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05029_));
 sky130_fd_sc_hd__nand2_1 _11231_ (.A(_04987_),
    .B(_05029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05030_));
 sky130_fd_sc_hd__o22a_1 _11232_ (.A1(net42),
    .A2(_04773_),
    .B1(_05024_),
    .B2(_05030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00130_));
 sky130_fd_sc_hd__mux4_1 _11233_ (.A0(\fifo_inst.mem.rMemory[8][21] ),
    .A1(\fifo_inst.mem.rMemory[9][21] ),
    .A2(\fifo_inst.mem.rMemory[10][21] ),
    .A3(\fifo_inst.mem.rMemory[11][21] ),
    .S0(_05008_),
    .S1(_05009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05031_));
 sky130_fd_sc_hd__mux4_1 _11234_ (.A0(\fifo_inst.mem.rMemory[12][21] ),
    .A1(\fifo_inst.mem.rMemory[13][21] ),
    .A2(\fifo_inst.mem.rMemory[14][21] ),
    .A3(\fifo_inst.mem.rMemory[15][21] ),
    .S0(_04807_),
    .S1(_04809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05032_));
 sky130_fd_sc_hd__or2b_1 _11235_ (.A(_05032_),
    .B_N(_04776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05033_));
 sky130_fd_sc_hd__o211a_1 _11236_ (.A1(_05007_),
    .A2(_05031_),
    .B1(_05033_),
    .C1(_05023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05034_));
 sky130_fd_sc_hd__mux4_1 _11237_ (.A0(\fifo_inst.mem.rMemory[4][21] ),
    .A1(\fifo_inst.mem.rMemory[5][21] ),
    .A2(\fifo_inst.mem.rMemory[6][21] ),
    .A3(\fifo_inst.mem.rMemory[7][21] ),
    .S0(_04988_),
    .S1(_04989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05035_));
 sky130_fd_sc_hd__inv_2 _11238_ (.A(_05035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05036_));
 sky130_fd_sc_hd__mux4_1 _11239_ (.A0(\fifo_inst.mem.rMemory[0][21] ),
    .A1(\fifo_inst.mem.rMemory[1][21] ),
    .A2(\fifo_inst.mem.rMemory[2][21] ),
    .A3(\fifo_inst.mem.rMemory[3][21] ),
    .S0(_04732_),
    .S1(_04736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05037_));
 sky130_fd_sc_hd__nor2_1 _11240_ (.A(_04992_),
    .B(_05037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05038_));
 sky130_fd_sc_hd__a211o_1 _11241_ (.A1(_04758_),
    .A2(_05036_),
    .B1(_05038_),
    .C1(_04747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05039_));
 sky130_fd_sc_hd__nand2_1 _11242_ (.A(_04987_),
    .B(_05039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05040_));
 sky130_fd_sc_hd__o22a_1 _11243_ (.A1(net43),
    .A2(_04773_),
    .B1(_05034_),
    .B2(_05040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00131_));
 sky130_fd_sc_hd__mux4_1 _11244_ (.A0(\fifo_inst.mem.rMemory[8][22] ),
    .A1(\fifo_inst.mem.rMemory[9][22] ),
    .A2(\fifo_inst.mem.rMemory[10][22] ),
    .A3(\fifo_inst.mem.rMemory[11][22] ),
    .S0(_05008_),
    .S1(_05009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05041_));
 sky130_fd_sc_hd__mux4_1 _11245_ (.A0(\fifo_inst.mem.rMemory[12][22] ),
    .A1(\fifo_inst.mem.rMemory[13][22] ),
    .A2(\fifo_inst.mem.rMemory[14][22] ),
    .A3(\fifo_inst.mem.rMemory[15][22] ),
    .S0(_04807_),
    .S1(_04809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05042_));
 sky130_fd_sc_hd__or2b_1 _11246_ (.A(_05042_),
    .B_N(_04776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05043_));
 sky130_fd_sc_hd__o211a_1 _11247_ (.A1(_05007_),
    .A2(_05041_),
    .B1(_05043_),
    .C1(_05023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05044_));
 sky130_fd_sc_hd__mux4_1 _11248_ (.A0(\fifo_inst.mem.rMemory[4][22] ),
    .A1(\fifo_inst.mem.rMemory[5][22] ),
    .A2(\fifo_inst.mem.rMemory[6][22] ),
    .A3(\fifo_inst.mem.rMemory[7][22] ),
    .S0(_04731_),
    .S1(_04760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05045_));
 sky130_fd_sc_hd__inv_2 _11249_ (.A(_05045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05046_));
 sky130_fd_sc_hd__mux4_1 _11250_ (.A0(\fifo_inst.mem.rMemory[0][22] ),
    .A1(\fifo_inst.mem.rMemory[1][22] ),
    .A2(\fifo_inst.mem.rMemory[2][22] ),
    .A3(\fifo_inst.mem.rMemory[3][22] ),
    .S0(_04732_),
    .S1(_04736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05047_));
 sky130_fd_sc_hd__nor2_1 _11251_ (.A(_04728_),
    .B(_05047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05048_));
 sky130_fd_sc_hd__a211o_1 _11252_ (.A1(_04758_),
    .A2(_05046_),
    .B1(_05048_),
    .C1(_04747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05049_));
 sky130_fd_sc_hd__nand2_1 _11253_ (.A(_04725_),
    .B(_05049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05050_));
 sky130_fd_sc_hd__o22a_1 _11254_ (.A1(net44),
    .A2(_04773_),
    .B1(_05044_),
    .B2(_05050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00132_));
 sky130_fd_sc_hd__mux4_1 _11255_ (.A0(\fifo_inst.mem.rMemory[8][23] ),
    .A1(\fifo_inst.mem.rMemory[9][23] ),
    .A2(\fifo_inst.mem.rMemory[10][23] ),
    .A3(\fifo_inst.mem.rMemory[11][23] ),
    .S0(_05008_),
    .S1(_05009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05051_));
 sky130_fd_sc_hd__mux4_1 _11256_ (.A0(\fifo_inst.mem.rMemory[12][23] ),
    .A1(\fifo_inst.mem.rMemory[13][23] ),
    .A2(\fifo_inst.mem.rMemory[14][23] ),
    .A3(\fifo_inst.mem.rMemory[15][23] ),
    .S0(_04807_),
    .S1(_04809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05052_));
 sky130_fd_sc_hd__or2b_1 _11257_ (.A(_05052_),
    .B_N(_04776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05053_));
 sky130_fd_sc_hd__o211a_1 _11258_ (.A1(_05007_),
    .A2(_05051_),
    .B1(_05053_),
    .C1(_05023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05054_));
 sky130_fd_sc_hd__mux4_1 _11259_ (.A0(\fifo_inst.mem.rMemory[4][23] ),
    .A1(\fifo_inst.mem.rMemory[5][23] ),
    .A2(\fifo_inst.mem.rMemory[6][23] ),
    .A3(\fifo_inst.mem.rMemory[7][23] ),
    .S0(_04731_),
    .S1(_04760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05055_));
 sky130_fd_sc_hd__inv_2 _11260_ (.A(_05055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05056_));
 sky130_fd_sc_hd__mux4_1 _11261_ (.A0(\fifo_inst.mem.rMemory[0][23] ),
    .A1(\fifo_inst.mem.rMemory[1][23] ),
    .A2(\fifo_inst.mem.rMemory[2][23] ),
    .A3(\fifo_inst.mem.rMemory[3][23] ),
    .S0(_04732_),
    .S1(_04736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05057_));
 sky130_fd_sc_hd__nor2_1 _11262_ (.A(_04728_),
    .B(_05057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05058_));
 sky130_fd_sc_hd__a211o_1 _11263_ (.A1(_04758_),
    .A2(_05056_),
    .B1(_05058_),
    .C1(_04747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05059_));
 sky130_fd_sc_hd__nand2_1 _11264_ (.A(_04725_),
    .B(_05059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05060_));
 sky130_fd_sc_hd__o22a_1 _11265_ (.A1(net45),
    .A2(_04773_),
    .B1(_05054_),
    .B2(_05060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00133_));
 sky130_fd_sc_hd__and2_1 _11266_ (.A(_02163_),
    .B(_02154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05061_));
 sky130_fd_sc_hd__clkbuf_1 _11267_ (.A(_05061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00134_));
 sky130_fd_sc_hd__and2_1 _11268_ (.A(_03194_),
    .B(_03185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05062_));
 sky130_fd_sc_hd__clkbuf_1 _11269_ (.A(_05062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00135_));
 sky130_fd_sc_hd__and2b_1 _11270_ (.A_N(_04138_),
    .B(_04135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05063_));
 sky130_fd_sc_hd__clkbuf_1 _11271_ (.A(_05063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00136_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11272_ (.A(\fifo_inst.WR_DATA[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05064_));
 sky130_fd_sc_hd__clkbuf_2 _11273_ (.A(\fifo_inst.mem.WR1_ADDR[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05065_));
 sky130_fd_sc_hd__inv_2 _11274_ (.A(\fifo_inst.rFull ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05066_));
 sky130_fd_sc_hd__o31ai_4 _11275_ (.A1(\shift_register[10] ),
    .A2(\shift_register[9] ),
    .A3(\shift_register[11] ),
    .B1(_05066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05067_));
 sky130_fd_sc_hd__or3b_4 _11276_ (.A(_05065_),
    .B(_05067_),
    .C_N(\fifo_inst.mem.WR1_ADDR[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05068_));
 sky130_fd_sc_hd__buf_2 _11277_ (.A(\fifo_inst.mem.WR1_ADDR[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05069_));
 sky130_fd_sc_hd__buf_2 _11278_ (.A(\fifo_inst.mem.WR1_ADDR[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05070_));
 sky130_fd_sc_hd__or2_4 _11279_ (.A(_05069_),
    .B(_05070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05071_));
 sky130_fd_sc_hd__nor2_8 _11280_ (.A(_05068_),
    .B(_05071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05072_));
 sky130_fd_sc_hd__clkbuf_2 _11281_ (.A(_05072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05073_));
 sky130_fd_sc_hd__buf_2 _11282_ (.A(_05073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05074_));
 sky130_fd_sc_hd__mux2_1 _11283_ (.A0(\fifo_inst.mem.rMemory[2][0] ),
    .A1(_05064_),
    .S(_05074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05075_));
 sky130_fd_sc_hd__clkbuf_1 _11284_ (.A(_05075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00137_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11285_ (.A(\fifo_inst.WR_DATA[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05076_));
 sky130_fd_sc_hd__mux2_1 _11286_ (.A0(\fifo_inst.mem.rMemory[2][1] ),
    .A1(_05076_),
    .S(_05074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05077_));
 sky130_fd_sc_hd__clkbuf_1 _11287_ (.A(_05077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00138_));
 sky130_fd_sc_hd__clkbuf_2 _11288_ (.A(\fifo_inst.WR_DATA[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05078_));
 sky130_fd_sc_hd__mux2_1 _11289_ (.A0(\fifo_inst.mem.rMemory[2][2] ),
    .A1(_05078_),
    .S(_05074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05079_));
 sky130_fd_sc_hd__clkbuf_1 _11290_ (.A(_05079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00139_));
 sky130_fd_sc_hd__clkbuf_2 _11291_ (.A(\fifo_inst.WR_DATA[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05080_));
 sky130_fd_sc_hd__mux2_1 _11292_ (.A0(\fifo_inst.mem.rMemory[2][3] ),
    .A1(_05080_),
    .S(_05074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05081_));
 sky130_fd_sc_hd__clkbuf_1 _11293_ (.A(_05081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00140_));
 sky130_fd_sc_hd__clkbuf_2 _11294_ (.A(\fifo_inst.WR_DATA[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05082_));
 sky130_fd_sc_hd__mux2_1 _11295_ (.A0(\fifo_inst.mem.rMemory[2][4] ),
    .A1(_05082_),
    .S(_05074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05083_));
 sky130_fd_sc_hd__clkbuf_1 _11296_ (.A(_05083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00141_));
 sky130_fd_sc_hd__buf_2 _11297_ (.A(\fifo_inst.WR_DATA[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05084_));
 sky130_fd_sc_hd__buf_2 _11298_ (.A(_05072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05085_));
 sky130_fd_sc_hd__mux2_1 _11299_ (.A0(\fifo_inst.mem.rMemory[2][5] ),
    .A1(_05084_),
    .S(_05085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05086_));
 sky130_fd_sc_hd__clkbuf_1 _11300_ (.A(_05086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00142_));
 sky130_fd_sc_hd__clkbuf_2 _11301_ (.A(\fifo_inst.WR_DATA[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05087_));
 sky130_fd_sc_hd__mux2_1 _11302_ (.A0(\fifo_inst.mem.rMemory[2][6] ),
    .A1(_05087_),
    .S(_05085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05088_));
 sky130_fd_sc_hd__clkbuf_1 _11303_ (.A(_05088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00143_));
 sky130_fd_sc_hd__buf_2 _11304_ (.A(\fifo_inst.WR_DATA[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05089_));
 sky130_fd_sc_hd__mux2_1 _11305_ (.A0(\fifo_inst.mem.rMemory[2][7] ),
    .A1(_05089_),
    .S(_05085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05090_));
 sky130_fd_sc_hd__clkbuf_1 _11306_ (.A(_05090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00144_));
 sky130_fd_sc_hd__buf_2 _11307_ (.A(\fifo_inst.WR_DATA[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05091_));
 sky130_fd_sc_hd__mux2_1 _11308_ (.A0(\fifo_inst.mem.rMemory[2][8] ),
    .A1(_05091_),
    .S(_05085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05092_));
 sky130_fd_sc_hd__clkbuf_1 _11309_ (.A(_05092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00145_));
 sky130_fd_sc_hd__clkbuf_2 _11310_ (.A(\fifo_inst.WR_DATA[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05093_));
 sky130_fd_sc_hd__mux2_1 _11311_ (.A0(\fifo_inst.mem.rMemory[2][9] ),
    .A1(_05093_),
    .S(_05085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05094_));
 sky130_fd_sc_hd__clkbuf_1 _11312_ (.A(_05094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00146_));
 sky130_fd_sc_hd__clkbuf_2 _11313_ (.A(\fifo_inst.WR_DATA[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05095_));
 sky130_fd_sc_hd__buf_2 _11314_ (.A(_05072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05096_));
 sky130_fd_sc_hd__mux2_1 _11315_ (.A0(\fifo_inst.mem.rMemory[2][10] ),
    .A1(_05095_),
    .S(_05096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05097_));
 sky130_fd_sc_hd__clkbuf_1 _11316_ (.A(_05097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00147_));
 sky130_fd_sc_hd__clkbuf_2 _11317_ (.A(\fifo_inst.WR_DATA[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05098_));
 sky130_fd_sc_hd__mux2_1 _11318_ (.A0(\fifo_inst.mem.rMemory[2][11] ),
    .A1(_05098_),
    .S(_05096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05099_));
 sky130_fd_sc_hd__clkbuf_1 _11319_ (.A(_05099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00148_));
 sky130_fd_sc_hd__clkbuf_2 _11320_ (.A(\fifo_inst.WR_DATA[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05100_));
 sky130_fd_sc_hd__mux2_1 _11321_ (.A0(\fifo_inst.mem.rMemory[2][12] ),
    .A1(_05100_),
    .S(_05096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05101_));
 sky130_fd_sc_hd__clkbuf_1 _11322_ (.A(_05101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00149_));
 sky130_fd_sc_hd__buf_2 _11323_ (.A(\fifo_inst.WR_DATA[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05102_));
 sky130_fd_sc_hd__mux2_1 _11324_ (.A0(\fifo_inst.mem.rMemory[2][13] ),
    .A1(_05102_),
    .S(_05096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05103_));
 sky130_fd_sc_hd__clkbuf_1 _11325_ (.A(_05103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00150_));
 sky130_fd_sc_hd__buf_2 _11326_ (.A(\fifo_inst.WR_DATA[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05104_));
 sky130_fd_sc_hd__mux2_1 _11327_ (.A0(\fifo_inst.mem.rMemory[2][14] ),
    .A1(_05104_),
    .S(_05096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05105_));
 sky130_fd_sc_hd__clkbuf_1 _11328_ (.A(_05105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00151_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11329_ (.A(\fifo_inst.WR_DATA[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05106_));
 sky130_fd_sc_hd__buf_2 _11330_ (.A(_05072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05107_));
 sky130_fd_sc_hd__mux2_1 _11331_ (.A0(\fifo_inst.mem.rMemory[2][15] ),
    .A1(_05106_),
    .S(_05107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05108_));
 sky130_fd_sc_hd__clkbuf_1 _11332_ (.A(_05108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00152_));
 sky130_fd_sc_hd__nor2_1 _11333_ (.A(\sa_inst.cols_l2a:3.l2a_i._23_ ),
    .B(\sa_inst.cols_l2a:3.l2a_i._27_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05109_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11334_ (.A(_05109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05110_));
 sky130_fd_sc_hd__o21ai_1 _11335_ (.A1(\sa_inst.cols_l2a:3.l2a_i._09_[0] ),
    .A2(\sa_inst.cols_l2a:3.l2a_i._15_ ),
    .B1(_05110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05111_));
 sky130_fd_sc_hd__a21oi_4 _11336_ (.A1(\sa_inst.cols_l2a:3.l2a_i._09_[0] ),
    .A2(\sa_inst.cols_l2a:3.l2a_i._15_ ),
    .B1(_05111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05112_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11337_ (.A(_05112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05113_));
 sky130_fd_sc_hd__mux2_1 _11338_ (.A0(\fifo_inst.mem.rMemory[2][16] ),
    .A1(_05113_),
    .S(_05107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05114_));
 sky130_fd_sc_hd__clkbuf_1 _11339_ (.A(_05114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00153_));
 sky130_fd_sc_hd__and3_1 _11340_ (.A(\sa_inst.cols_l2a:3.l2a_i._09_[0] ),
    .B(\sa_inst.cols_l2a:3.l2a_i._15_ ),
    .C(\sa_inst.cols_l2a:3.l2a_i._09_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05115_));
 sky130_fd_sc_hd__a21o_1 _11341_ (.A1(\sa_inst.cols_l2a:3.l2a_i._09_[0] ),
    .A2(\sa_inst.cols_l2a:3.l2a_i._15_ ),
    .B1(\sa_inst.cols_l2a:3.l2a_i._09_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05116_));
 sky130_fd_sc_hd__and3b_4 _11342_ (.A_N(_05115_),
    .B(_05110_),
    .C(_05116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05117_));
 sky130_fd_sc_hd__clkbuf_2 _11343_ (.A(_05117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05118_));
 sky130_fd_sc_hd__mux2_1 _11344_ (.A0(\fifo_inst.mem.rMemory[2][17] ),
    .A1(_05118_),
    .S(_05107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05119_));
 sky130_fd_sc_hd__clkbuf_1 _11345_ (.A(_05119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00154_));
 sky130_fd_sc_hd__o21ai_1 _11346_ (.A1(\sa_inst.cols_l2a:3.l2a_i._09_[2] ),
    .A2(_05115_),
    .B1(_05110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05120_));
 sky130_fd_sc_hd__a21oi_4 _11347_ (.A1(\sa_inst.cols_l2a:3.l2a_i._09_[2] ),
    .A2(_05115_),
    .B1(_05120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05121_));
 sky130_fd_sc_hd__clkbuf_2 _11348_ (.A(_05121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05122_));
 sky130_fd_sc_hd__mux2_1 _11349_ (.A0(\fifo_inst.mem.rMemory[2][18] ),
    .A1(_05122_),
    .S(_05107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05123_));
 sky130_fd_sc_hd__clkbuf_1 _11350_ (.A(_05123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00155_));
 sky130_fd_sc_hd__and3_2 _11351_ (.A(\sa_inst.cols_l2a:3.l2a_i._09_[2] ),
    .B(\sa_inst.cols_l2a:3.l2a_i._09_[3] ),
    .C(_05115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05124_));
 sky130_fd_sc_hd__a21o_1 _11352_ (.A1(\sa_inst.cols_l2a:3.l2a_i._09_[2] ),
    .A2(_05115_),
    .B1(\sa_inst.cols_l2a:3.l2a_i._09_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05125_));
 sky130_fd_sc_hd__and3b_4 _11353_ (.A_N(_05124_),
    .B(_05110_),
    .C(_05125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05126_));
 sky130_fd_sc_hd__clkbuf_2 _11354_ (.A(_05126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05127_));
 sky130_fd_sc_hd__mux2_1 _11355_ (.A0(\fifo_inst.mem.rMemory[2][19] ),
    .A1(_05127_),
    .S(_05107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05128_));
 sky130_fd_sc_hd__clkbuf_1 _11356_ (.A(_05128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00156_));
 sky130_fd_sc_hd__o21ai_1 _11357_ (.A1(\sa_inst.cols_l2a:3.l2a_i._09_[4] ),
    .A2(_05124_),
    .B1(_05110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05129_));
 sky130_fd_sc_hd__a21oi_4 _11358_ (.A1(\sa_inst.cols_l2a:3.l2a_i._09_[4] ),
    .A2(_05124_),
    .B1(_05129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05130_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11359_ (.A(_05130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05131_));
 sky130_fd_sc_hd__mux2_1 _11360_ (.A0(\fifo_inst.mem.rMemory[2][20] ),
    .A1(_05131_),
    .S(_05073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05132_));
 sky130_fd_sc_hd__clkbuf_1 _11361_ (.A(_05132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00157_));
 sky130_fd_sc_hd__and3_1 _11362_ (.A(\sa_inst.cols_l2a:3.l2a_i._09_[4] ),
    .B(\sa_inst.cols_l2a:3.l2a_i._09_[5] ),
    .C(_05124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05133_));
 sky130_fd_sc_hd__a21o_1 _11363_ (.A1(\sa_inst.cols_l2a:3.l2a_i._09_[4] ),
    .A2(_05124_),
    .B1(\sa_inst.cols_l2a:3.l2a_i._09_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05134_));
 sky130_fd_sc_hd__and3b_4 _11364_ (.A_N(_05133_),
    .B(_05109_),
    .C(_05134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05135_));
 sky130_fd_sc_hd__clkbuf_2 _11365_ (.A(_05135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05136_));
 sky130_fd_sc_hd__mux2_1 _11366_ (.A0(\fifo_inst.mem.rMemory[2][21] ),
    .A1(_05136_),
    .S(_05073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05137_));
 sky130_fd_sc_hd__clkbuf_1 _11367_ (.A(_05137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00158_));
 sky130_fd_sc_hd__a21boi_1 _11368_ (.A1(\sa_inst.cols_l2a:3.l2a_i._09_[6] ),
    .A2(_05133_),
    .B1_N(_05109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05138_));
 sky130_fd_sc_hd__o21a_4 _11369_ (.A1(\sa_inst.cols_l2a:3.l2a_i._09_[6] ),
    .A2(_05133_),
    .B1(_05138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05139_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11370_ (.A(_05139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05140_));
 sky130_fd_sc_hd__mux2_1 _11371_ (.A0(\fifo_inst.mem.rMemory[2][22] ),
    .A1(_05140_),
    .S(_05073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05141_));
 sky130_fd_sc_hd__clkbuf_1 _11372_ (.A(_05141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00159_));
 sky130_fd_sc_hd__inv_2 _11373_ (.A(\sa_inst.cols_l2a:3.l2a_i._27_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05142_));
 sky130_fd_sc_hd__a21o_4 _11374_ (.A1(_05142_),
    .A2(\sa_inst.cols_l2a:3.l2a_i._55_ ),
    .B1(\sa_inst.cols_l2a:3.l2a_i._23_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05143_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11375_ (.A(_05143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05144_));
 sky130_fd_sc_hd__mux2_1 _11376_ (.A0(\fifo_inst.mem.rMemory[2][23] ),
    .A1(_05144_),
    .S(_05073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05145_));
 sky130_fd_sc_hd__clkbuf_1 _11377_ (.A(_05145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00160_));
 sky130_fd_sc_hd__and2_1 _11378_ (.A(\sa_inst._12_[67] ),
    .B(_00722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05146_));
 sky130_fd_sc_hd__clkbuf_1 _11379_ (.A(_05146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00161_));
 sky130_fd_sc_hd__and2_1 _11380_ (.A(\sa_inst._12_[68] ),
    .B(_00722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05147_));
 sky130_fd_sc_hd__clkbuf_1 _11381_ (.A(_05147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00162_));
 sky130_fd_sc_hd__and2_1 _11382_ (.A(\sa_inst._12_[69] ),
    .B(_00722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05148_));
 sky130_fd_sc_hd__clkbuf_1 _11383_ (.A(_05148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00163_));
 sky130_fd_sc_hd__clkbuf_2 _11384_ (.A(_00721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05149_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11385_ (.A(_05149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05150_));
 sky130_fd_sc_hd__and2_1 _11386_ (.A(\sa_inst._12_[70] ),
    .B(_05150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05151_));
 sky130_fd_sc_hd__clkbuf_1 _11387_ (.A(_05151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00164_));
 sky130_fd_sc_hd__and2_1 _11388_ (.A(\sa_inst._12_[71] ),
    .B(_05150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05152_));
 sky130_fd_sc_hd__clkbuf_1 _11389_ (.A(_05152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00165_));
 sky130_fd_sc_hd__and2_1 _11390_ (.A(\sa_inst._12_[72] ),
    .B(_05150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05153_));
 sky130_fd_sc_hd__clkbuf_1 _11391_ (.A(_05153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00166_));
 sky130_fd_sc_hd__and2_1 _11392_ (.A(\sa_inst._12_[73] ),
    .B(_05150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05154_));
 sky130_fd_sc_hd__clkbuf_1 _11393_ (.A(_05154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00167_));
 sky130_fd_sc_hd__and2_1 _11394_ (.A(\sa_inst._12_[74] ),
    .B(_05150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05155_));
 sky130_fd_sc_hd__clkbuf_1 _11395_ (.A(_05155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00168_));
 sky130_fd_sc_hd__clkbuf_1 _11396_ (.A(_05149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05156_));
 sky130_fd_sc_hd__and2_1 _11397_ (.A(\sa_inst._12_[75] ),
    .B(_05156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05157_));
 sky130_fd_sc_hd__clkbuf_1 _11398_ (.A(_05157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00169_));
 sky130_fd_sc_hd__and2_1 _11399_ (.A(\sa_inst._12_[76] ),
    .B(_05156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05158_));
 sky130_fd_sc_hd__clkbuf_1 _11400_ (.A(_05158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00170_));
 sky130_fd_sc_hd__and2_1 _11401_ (.A(\sa_inst._12_[77] ),
    .B(_05156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05159_));
 sky130_fd_sc_hd__clkbuf_1 _11402_ (.A(_05159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00171_));
 sky130_fd_sc_hd__and2_1 _11403_ (.A(\sa_inst._12_[78] ),
    .B(_05156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05160_));
 sky130_fd_sc_hd__clkbuf_1 _11404_ (.A(_05160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00172_));
 sky130_fd_sc_hd__and2_1 _11405_ (.A(\sa_inst._12_[79] ),
    .B(_05156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05161_));
 sky130_fd_sc_hd__clkbuf_1 _11406_ (.A(_05161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00173_));
 sky130_fd_sc_hd__clkbuf_1 _11407_ (.A(_00721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05162_));
 sky130_fd_sc_hd__and2_1 _11408_ (.A(\sa_inst._12_[80] ),
    .B(_05162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05163_));
 sky130_fd_sc_hd__clkbuf_1 _11409_ (.A(_05163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00174_));
 sky130_fd_sc_hd__and2_1 _11410_ (.A(\sa_inst._12_[81] ),
    .B(_05162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05164_));
 sky130_fd_sc_hd__clkbuf_1 _11411_ (.A(_05164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00175_));
 sky130_fd_sc_hd__and2_1 _11412_ (.A(\sa_inst._12_[82] ),
    .B(_05162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05165_));
 sky130_fd_sc_hd__clkbuf_1 _11413_ (.A(_05165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00176_));
 sky130_fd_sc_hd__and2_1 _11414_ (.A(\sa_inst._12_[83] ),
    .B(_05162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05166_));
 sky130_fd_sc_hd__clkbuf_1 _11415_ (.A(_05166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00177_));
 sky130_fd_sc_hd__and2_1 _11416_ (.A(\sa_inst._12_[84] ),
    .B(_05162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05167_));
 sky130_fd_sc_hd__clkbuf_1 _11417_ (.A(_05167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00178_));
 sky130_fd_sc_hd__clkbuf_1 _11418_ (.A(_00721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05168_));
 sky130_fd_sc_hd__and2_1 _11419_ (.A(\sa_inst._12_[85] ),
    .B(_05168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05169_));
 sky130_fd_sc_hd__clkbuf_1 _11420_ (.A(_05169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00179_));
 sky130_fd_sc_hd__and2_1 _11421_ (.A(\sa_inst._12_[86] ),
    .B(_05168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05170_));
 sky130_fd_sc_hd__clkbuf_1 _11422_ (.A(_05170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00180_));
 sky130_fd_sc_hd__and2_1 _11423_ (.A(\sa_inst._12_[87] ),
    .B(_05168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05171_));
 sky130_fd_sc_hd__clkbuf_1 _11424_ (.A(_05171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00181_));
 sky130_fd_sc_hd__and2_1 _11425_ (.A(\sa_inst._12_[88] ),
    .B(_05168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05172_));
 sky130_fd_sc_hd__clkbuf_1 _11426_ (.A(_05172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00182_));
 sky130_fd_sc_hd__and2_1 _11427_ (.A(\sa_inst._12_[89] ),
    .B(_05168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05173_));
 sky130_fd_sc_hd__clkbuf_1 _11428_ (.A(_05173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00183_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11429_ (.A(_00721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05174_));
 sky130_fd_sc_hd__and2_1 _11430_ (.A(\sa_inst._12_[90] ),
    .B(_05174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05175_));
 sky130_fd_sc_hd__clkbuf_1 _11431_ (.A(_05175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00184_));
 sky130_fd_sc_hd__and2_1 _11432_ (.A(\sa_inst._12_[91] ),
    .B(_05174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05176_));
 sky130_fd_sc_hd__clkbuf_1 _11433_ (.A(_05176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00185_));
 sky130_fd_sc_hd__and2_1 _11434_ (.A(\sa_inst._12_[92] ),
    .B(_05174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05177_));
 sky130_fd_sc_hd__clkbuf_1 _11435_ (.A(_05177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00186_));
 sky130_fd_sc_hd__and2_1 _11436_ (.A(\sa_inst._12_[93] ),
    .B(_05174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05178_));
 sky130_fd_sc_hd__clkbuf_1 _11437_ (.A(_05178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00187_));
 sky130_fd_sc_hd__and2_1 _11438_ (.A(\sa_inst._12_[94] ),
    .B(_05174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05179_));
 sky130_fd_sc_hd__clkbuf_1 _11439_ (.A(_05179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00188_));
 sky130_fd_sc_hd__and2_1 _11440_ (.A(\sa_inst._12_[95] ),
    .B(_05149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05180_));
 sky130_fd_sc_hd__clkbuf_1 _11441_ (.A(_05180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00189_));
 sky130_fd_sc_hd__and2_1 _11442_ (.A(\sa_inst._12_[96] ),
    .B(_05149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05181_));
 sky130_fd_sc_hd__clkbuf_1 _11443_ (.A(_05181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00190_));
 sky130_fd_sc_hd__and2_1 _11444_ (.A(\sa_inst._12_[97] ),
    .B(_05149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05182_));
 sky130_fd_sc_hd__clkbuf_1 _11445_ (.A(_05182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00191_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11446_ (.A(\fifo_inst.WR_DATA[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05183_));
 sky130_fd_sc_hd__nand2_8 _11447_ (.A(_05069_),
    .B(_05070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05184_));
 sky130_fd_sc_hd__nor2_8 _11448_ (.A(_05068_),
    .B(_05184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05185_));
 sky130_fd_sc_hd__buf_2 _11449_ (.A(_05185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05186_));
 sky130_fd_sc_hd__buf_2 _11450_ (.A(_05186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05187_));
 sky130_fd_sc_hd__mux2_1 _11451_ (.A0(\fifo_inst.mem.rMemory[14][0] ),
    .A1(_05183_),
    .S(_05187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05188_));
 sky130_fd_sc_hd__clkbuf_1 _11452_ (.A(_05188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00192_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11453_ (.A(\fifo_inst.WR_DATA[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05189_));
 sky130_fd_sc_hd__mux2_1 _11454_ (.A0(\fifo_inst.mem.rMemory[14][1] ),
    .A1(_05189_),
    .S(_05187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05190_));
 sky130_fd_sc_hd__clkbuf_1 _11455_ (.A(_05190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00193_));
 sky130_fd_sc_hd__clkbuf_2 _11456_ (.A(\fifo_inst.WR_DATA[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05191_));
 sky130_fd_sc_hd__mux2_1 _11457_ (.A0(\fifo_inst.mem.rMemory[14][2] ),
    .A1(_05191_),
    .S(_05187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05192_));
 sky130_fd_sc_hd__clkbuf_1 _11458_ (.A(_05192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00194_));
 sky130_fd_sc_hd__clkbuf_2 _11459_ (.A(\fifo_inst.WR_DATA[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05193_));
 sky130_fd_sc_hd__mux2_1 _11460_ (.A0(\fifo_inst.mem.rMemory[14][3] ),
    .A1(_05193_),
    .S(_05187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05194_));
 sky130_fd_sc_hd__clkbuf_1 _11461_ (.A(_05194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00195_));
 sky130_fd_sc_hd__clkbuf_2 _11462_ (.A(\fifo_inst.WR_DATA[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05195_));
 sky130_fd_sc_hd__mux2_1 _11463_ (.A0(\fifo_inst.mem.rMemory[14][4] ),
    .A1(_05195_),
    .S(_05187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05196_));
 sky130_fd_sc_hd__clkbuf_1 _11464_ (.A(_05196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00196_));
 sky130_fd_sc_hd__clkbuf_2 _11465_ (.A(\fifo_inst.WR_DATA[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05197_));
 sky130_fd_sc_hd__buf_2 _11466_ (.A(_05185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05198_));
 sky130_fd_sc_hd__mux2_1 _11467_ (.A0(\fifo_inst.mem.rMemory[14][5] ),
    .A1(_05197_),
    .S(_05198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05199_));
 sky130_fd_sc_hd__clkbuf_1 _11468_ (.A(_05199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00197_));
 sky130_fd_sc_hd__clkbuf_2 _11469_ (.A(\fifo_inst.WR_DATA[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05200_));
 sky130_fd_sc_hd__mux2_1 _11470_ (.A0(\fifo_inst.mem.rMemory[14][6] ),
    .A1(_05200_),
    .S(_05198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05201_));
 sky130_fd_sc_hd__clkbuf_1 _11471_ (.A(_05201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00198_));
 sky130_fd_sc_hd__buf_2 _11472_ (.A(\fifo_inst.WR_DATA[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05202_));
 sky130_fd_sc_hd__mux2_1 _11473_ (.A0(\fifo_inst.mem.rMemory[14][7] ),
    .A1(_05202_),
    .S(_05198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05203_));
 sky130_fd_sc_hd__clkbuf_1 _11474_ (.A(_05203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00199_));
 sky130_fd_sc_hd__clkbuf_2 _11475_ (.A(\fifo_inst.WR_DATA[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05204_));
 sky130_fd_sc_hd__mux2_1 _11476_ (.A0(\fifo_inst.mem.rMemory[14][8] ),
    .A1(_05204_),
    .S(_05198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05205_));
 sky130_fd_sc_hd__clkbuf_1 _11477_ (.A(_05205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00200_));
 sky130_fd_sc_hd__clkbuf_2 _11478_ (.A(\fifo_inst.WR_DATA[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05206_));
 sky130_fd_sc_hd__mux2_1 _11479_ (.A0(\fifo_inst.mem.rMemory[14][9] ),
    .A1(_05206_),
    .S(_05198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05207_));
 sky130_fd_sc_hd__clkbuf_1 _11480_ (.A(_05207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00201_));
 sky130_fd_sc_hd__clkbuf_2 _11481_ (.A(\fifo_inst.WR_DATA[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05208_));
 sky130_fd_sc_hd__buf_2 _11482_ (.A(_05185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05209_));
 sky130_fd_sc_hd__mux2_1 _11483_ (.A0(\fifo_inst.mem.rMemory[14][10] ),
    .A1(_05208_),
    .S(_05209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05210_));
 sky130_fd_sc_hd__clkbuf_1 _11484_ (.A(_05210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00202_));
 sky130_fd_sc_hd__clkbuf_2 _11485_ (.A(\fifo_inst.WR_DATA[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05211_));
 sky130_fd_sc_hd__mux2_1 _11486_ (.A0(\fifo_inst.mem.rMemory[14][11] ),
    .A1(_05211_),
    .S(_05209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05212_));
 sky130_fd_sc_hd__clkbuf_1 _11487_ (.A(_05212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00203_));
 sky130_fd_sc_hd__clkbuf_2 _11488_ (.A(\fifo_inst.WR_DATA[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05213_));
 sky130_fd_sc_hd__mux2_1 _11489_ (.A0(\fifo_inst.mem.rMemory[14][12] ),
    .A1(_05213_),
    .S(_05209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05214_));
 sky130_fd_sc_hd__clkbuf_1 _11490_ (.A(_05214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00204_));
 sky130_fd_sc_hd__buf_2 _11491_ (.A(\fifo_inst.WR_DATA[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05215_));
 sky130_fd_sc_hd__mux2_1 _11492_ (.A0(\fifo_inst.mem.rMemory[14][13] ),
    .A1(_05215_),
    .S(_05209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05216_));
 sky130_fd_sc_hd__clkbuf_1 _11493_ (.A(_05216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00205_));
 sky130_fd_sc_hd__buf_2 _11494_ (.A(\fifo_inst.WR_DATA[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05217_));
 sky130_fd_sc_hd__mux2_1 _11495_ (.A0(\fifo_inst.mem.rMemory[14][14] ),
    .A1(_05217_),
    .S(_05209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05218_));
 sky130_fd_sc_hd__clkbuf_1 _11496_ (.A(_05218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00206_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11497_ (.A(\fifo_inst.WR_DATA[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05219_));
 sky130_fd_sc_hd__buf_2 _11498_ (.A(_05185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05220_));
 sky130_fd_sc_hd__mux2_1 _11499_ (.A0(\fifo_inst.mem.rMemory[14][15] ),
    .A1(_05219_),
    .S(_05220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05221_));
 sky130_fd_sc_hd__clkbuf_1 _11500_ (.A(_05221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00207_));
 sky130_fd_sc_hd__clkbuf_2 _11501_ (.A(_05112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05222_));
 sky130_fd_sc_hd__mux2_1 _11502_ (.A0(\fifo_inst.mem.rMemory[14][16] ),
    .A1(_05222_),
    .S(_05220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05223_));
 sky130_fd_sc_hd__clkbuf_1 _11503_ (.A(_05223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00208_));
 sky130_fd_sc_hd__clkbuf_2 _11504_ (.A(_05117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05224_));
 sky130_fd_sc_hd__mux2_1 _11505_ (.A0(\fifo_inst.mem.rMemory[14][17] ),
    .A1(_05224_),
    .S(_05220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05225_));
 sky130_fd_sc_hd__clkbuf_1 _11506_ (.A(_05225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00209_));
 sky130_fd_sc_hd__clkbuf_2 _11507_ (.A(_05121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05226_));
 sky130_fd_sc_hd__mux2_1 _11508_ (.A0(\fifo_inst.mem.rMemory[14][18] ),
    .A1(_05226_),
    .S(_05220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05227_));
 sky130_fd_sc_hd__clkbuf_1 _11509_ (.A(_05227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00210_));
 sky130_fd_sc_hd__clkbuf_2 _11510_ (.A(_05126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05228_));
 sky130_fd_sc_hd__mux2_1 _11511_ (.A0(\fifo_inst.mem.rMemory[14][19] ),
    .A1(_05228_),
    .S(_05220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05229_));
 sky130_fd_sc_hd__clkbuf_1 _11512_ (.A(_05229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00211_));
 sky130_fd_sc_hd__clkbuf_2 _11513_ (.A(_05130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05230_));
 sky130_fd_sc_hd__mux2_1 _11514_ (.A0(\fifo_inst.mem.rMemory[14][20] ),
    .A1(_05230_),
    .S(_05186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05231_));
 sky130_fd_sc_hd__clkbuf_1 _11515_ (.A(_05231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00212_));
 sky130_fd_sc_hd__clkbuf_2 _11516_ (.A(_05135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05232_));
 sky130_fd_sc_hd__mux2_1 _11517_ (.A0(\fifo_inst.mem.rMemory[14][21] ),
    .A1(_05232_),
    .S(_05186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05233_));
 sky130_fd_sc_hd__clkbuf_1 _11518_ (.A(_05233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00213_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11519_ (.A(_05139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05234_));
 sky130_fd_sc_hd__mux2_1 _11520_ (.A0(\fifo_inst.mem.rMemory[14][22] ),
    .A1(_05234_),
    .S(_05186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05235_));
 sky130_fd_sc_hd__clkbuf_1 _11521_ (.A(_05235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00214_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11522_ (.A(_05143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05236_));
 sky130_fd_sc_hd__mux2_1 _11523_ (.A0(\fifo_inst.mem.rMemory[14][23] ),
    .A1(_05236_),
    .S(_05186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05237_));
 sky130_fd_sc_hd__clkbuf_1 _11524_ (.A(_05237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00215_));
 sky130_fd_sc_hd__and2_1 _11525_ (.A(\sa_inst._12_[34] ),
    .B(_00762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05238_));
 sky130_fd_sc_hd__clkbuf_1 _11526_ (.A(_05238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00216_));
 sky130_fd_sc_hd__and2_1 _11527_ (.A(\sa_inst._12_[35] ),
    .B(_00762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05239_));
 sky130_fd_sc_hd__clkbuf_1 _11528_ (.A(_05239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00217_));
 sky130_fd_sc_hd__and2_1 _11529_ (.A(\sa_inst._12_[36] ),
    .B(_00762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05240_));
 sky130_fd_sc_hd__clkbuf_1 _11530_ (.A(_05240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00218_));
 sky130_fd_sc_hd__clkbuf_2 _11531_ (.A(_00761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05241_));
 sky130_fd_sc_hd__clkbuf_1 _11532_ (.A(_05241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05242_));
 sky130_fd_sc_hd__and2_1 _11533_ (.A(\sa_inst._12_[37] ),
    .B(_05242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05243_));
 sky130_fd_sc_hd__clkbuf_1 _11534_ (.A(_05243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00219_));
 sky130_fd_sc_hd__and2_1 _11535_ (.A(\sa_inst._12_[38] ),
    .B(_05242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05244_));
 sky130_fd_sc_hd__clkbuf_1 _11536_ (.A(_05244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00220_));
 sky130_fd_sc_hd__and2_1 _11537_ (.A(\sa_inst._12_[39] ),
    .B(_05242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05245_));
 sky130_fd_sc_hd__clkbuf_1 _11538_ (.A(_05245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00221_));
 sky130_fd_sc_hd__and2_1 _11539_ (.A(\sa_inst._12_[40] ),
    .B(_05242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05246_));
 sky130_fd_sc_hd__clkbuf_1 _11540_ (.A(_05246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00222_));
 sky130_fd_sc_hd__and2_1 _11541_ (.A(\sa_inst._12_[41] ),
    .B(_05242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05247_));
 sky130_fd_sc_hd__clkbuf_1 _11542_ (.A(_05247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00223_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11543_ (.A(_05241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05248_));
 sky130_fd_sc_hd__and2_1 _11544_ (.A(\sa_inst._12_[42] ),
    .B(_05248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05249_));
 sky130_fd_sc_hd__clkbuf_1 _11545_ (.A(_05249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00224_));
 sky130_fd_sc_hd__and2_1 _11546_ (.A(\sa_inst._12_[43] ),
    .B(_05248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05250_));
 sky130_fd_sc_hd__clkbuf_1 _11547_ (.A(_05250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00225_));
 sky130_fd_sc_hd__and2_1 _11548_ (.A(\sa_inst._12_[44] ),
    .B(_05248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05251_));
 sky130_fd_sc_hd__clkbuf_1 _11549_ (.A(_05251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00226_));
 sky130_fd_sc_hd__and2_1 _11550_ (.A(\sa_inst._12_[45] ),
    .B(_05248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05252_));
 sky130_fd_sc_hd__clkbuf_1 _11551_ (.A(_05252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00227_));
 sky130_fd_sc_hd__and2_1 _11552_ (.A(\sa_inst._12_[46] ),
    .B(_05248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05253_));
 sky130_fd_sc_hd__clkbuf_1 _11553_ (.A(_05253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00228_));
 sky130_fd_sc_hd__clkbuf_1 _11554_ (.A(_00761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05254_));
 sky130_fd_sc_hd__and2_1 _11555_ (.A(\sa_inst._12_[47] ),
    .B(_05254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05255_));
 sky130_fd_sc_hd__clkbuf_1 _11556_ (.A(_05255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00229_));
 sky130_fd_sc_hd__and2_1 _11557_ (.A(\sa_inst._12_[48] ),
    .B(_05254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05256_));
 sky130_fd_sc_hd__clkbuf_1 _11558_ (.A(_05256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00230_));
 sky130_fd_sc_hd__and2_1 _11559_ (.A(\sa_inst._12_[49] ),
    .B(_05254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05257_));
 sky130_fd_sc_hd__clkbuf_1 _11560_ (.A(_05257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00231_));
 sky130_fd_sc_hd__and2_1 _11561_ (.A(\sa_inst._12_[50] ),
    .B(_05254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05258_));
 sky130_fd_sc_hd__clkbuf_1 _11562_ (.A(_05258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00232_));
 sky130_fd_sc_hd__and2_1 _11563_ (.A(\sa_inst._12_[51] ),
    .B(_05254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05259_));
 sky130_fd_sc_hd__clkbuf_1 _11564_ (.A(_05259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00233_));
 sky130_fd_sc_hd__clkbuf_1 _11565_ (.A(_00761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05260_));
 sky130_fd_sc_hd__and2_1 _11566_ (.A(\sa_inst._12_[52] ),
    .B(_05260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05261_));
 sky130_fd_sc_hd__clkbuf_1 _11567_ (.A(_05261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00234_));
 sky130_fd_sc_hd__and2_1 _11568_ (.A(\sa_inst._12_[53] ),
    .B(_05260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05262_));
 sky130_fd_sc_hd__clkbuf_1 _11569_ (.A(_05262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00235_));
 sky130_fd_sc_hd__and2_1 _11570_ (.A(\sa_inst._12_[54] ),
    .B(_05260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05263_));
 sky130_fd_sc_hd__clkbuf_1 _11571_ (.A(_05263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00236_));
 sky130_fd_sc_hd__and2_1 _11572_ (.A(\sa_inst._12_[55] ),
    .B(_05260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05264_));
 sky130_fd_sc_hd__clkbuf_1 _11573_ (.A(_05264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00237_));
 sky130_fd_sc_hd__and2_1 _11574_ (.A(\sa_inst._12_[56] ),
    .B(_05260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05265_));
 sky130_fd_sc_hd__clkbuf_1 _11575_ (.A(_05265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00238_));
 sky130_fd_sc_hd__clkbuf_1 _11576_ (.A(_00761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05266_));
 sky130_fd_sc_hd__and2_1 _11577_ (.A(\sa_inst._12_[57] ),
    .B(_05266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05267_));
 sky130_fd_sc_hd__clkbuf_1 _11578_ (.A(_05267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00239_));
 sky130_fd_sc_hd__and2_1 _11579_ (.A(\sa_inst._12_[58] ),
    .B(_05266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05268_));
 sky130_fd_sc_hd__clkbuf_1 _11580_ (.A(_05268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00240_));
 sky130_fd_sc_hd__and2_1 _11581_ (.A(\sa_inst._12_[59] ),
    .B(_05266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05269_));
 sky130_fd_sc_hd__clkbuf_1 _11582_ (.A(_05269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00241_));
 sky130_fd_sc_hd__and2_1 _11583_ (.A(\sa_inst._12_[60] ),
    .B(_05266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05270_));
 sky130_fd_sc_hd__clkbuf_1 _11584_ (.A(_05270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00242_));
 sky130_fd_sc_hd__and2_1 _11585_ (.A(\sa_inst._12_[61] ),
    .B(_05266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05271_));
 sky130_fd_sc_hd__clkbuf_1 _11586_ (.A(_05271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00243_));
 sky130_fd_sc_hd__and2_1 _11587_ (.A(\sa_inst._12_[62] ),
    .B(_05241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05272_));
 sky130_fd_sc_hd__clkbuf_1 _11588_ (.A(_05272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00244_));
 sky130_fd_sc_hd__and2_1 _11589_ (.A(\sa_inst._12_[63] ),
    .B(_05241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05273_));
 sky130_fd_sc_hd__clkbuf_1 _11590_ (.A(_05273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00245_));
 sky130_fd_sc_hd__and2_1 _11591_ (.A(\sa_inst._12_[64] ),
    .B(_05241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05274_));
 sky130_fd_sc_hd__clkbuf_1 _11592_ (.A(_05274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00246_));
 sky130_fd_sc_hd__and2_1 _11593_ (.A(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._03_ ),
    .B(_00858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05275_));
 sky130_fd_sc_hd__clkbuf_1 _11594_ (.A(_05275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00247_));
 sky130_fd_sc_hd__or4_1 _11595_ (.A(\sa_inst.cols_l2a:3.l2a_i._29_[0] ),
    .B(\sa_inst.cols_l2a:3.l2a_i._29_[1] ),
    .C(\sa_inst.cols_l2a:3.l2a_i._29_[3] ),
    .D(\sa_inst.cols_l2a:3.l2a_i._29_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05276_));
 sky130_fd_sc_hd__or4b_1 _11596_ (.A(\sa_inst.cols_l2a:3.l2a_i._29_[2] ),
    .B(\sa_inst.cols_l2a:3.l2a_i._29_[4] ),
    .C(_05276_),
    .D_N(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._55_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05277_));
 sky130_fd_sc_hd__inv_2 _11597_ (.A(_05277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00248_));
 sky130_fd_sc_hd__clkbuf_2 _11598_ (.A(\fifo_inst.mem.WR1_ADDR[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05278_));
 sky130_fd_sc_hd__inv_2 _11599_ (.A(_05065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05279_));
 sky130_fd_sc_hd__or3_4 _11600_ (.A(_05278_),
    .B(_05279_),
    .C(_05067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05280_));
 sky130_fd_sc_hd__nor2_8 _11601_ (.A(_05184_),
    .B(_05280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05281_));
 sky130_fd_sc_hd__buf_2 _11602_ (.A(_05281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05282_));
 sky130_fd_sc_hd__buf_2 _11603_ (.A(_05282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05283_));
 sky130_fd_sc_hd__mux2_1 _11604_ (.A0(\fifo_inst.mem.rMemory[13][0] ),
    .A1(_05183_),
    .S(_05283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05284_));
 sky130_fd_sc_hd__clkbuf_1 _11605_ (.A(_05284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _11606_ (.A0(\fifo_inst.mem.rMemory[13][1] ),
    .A1(_05189_),
    .S(_05283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05285_));
 sky130_fd_sc_hd__clkbuf_1 _11607_ (.A(_05285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _11608_ (.A0(\fifo_inst.mem.rMemory[13][2] ),
    .A1(_05191_),
    .S(_05283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05286_));
 sky130_fd_sc_hd__clkbuf_1 _11609_ (.A(_05286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _11610_ (.A0(\fifo_inst.mem.rMemory[13][3] ),
    .A1(_05193_),
    .S(_05283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05287_));
 sky130_fd_sc_hd__clkbuf_1 _11611_ (.A(_05287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _11612_ (.A0(\fifo_inst.mem.rMemory[13][4] ),
    .A1(_05195_),
    .S(_05283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05288_));
 sky130_fd_sc_hd__clkbuf_1 _11613_ (.A(_05288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00253_));
 sky130_fd_sc_hd__buf_2 _11614_ (.A(_05281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05289_));
 sky130_fd_sc_hd__mux2_1 _11615_ (.A0(\fifo_inst.mem.rMemory[13][5] ),
    .A1(_05197_),
    .S(_05289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05290_));
 sky130_fd_sc_hd__clkbuf_1 _11616_ (.A(_05290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _11617_ (.A0(\fifo_inst.mem.rMemory[13][6] ),
    .A1(_05200_),
    .S(_05289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05291_));
 sky130_fd_sc_hd__clkbuf_1 _11618_ (.A(_05291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _11619_ (.A0(\fifo_inst.mem.rMemory[13][7] ),
    .A1(_05202_),
    .S(_05289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05292_));
 sky130_fd_sc_hd__clkbuf_1 _11620_ (.A(_05292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _11621_ (.A0(\fifo_inst.mem.rMemory[13][8] ),
    .A1(_05204_),
    .S(_05289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05293_));
 sky130_fd_sc_hd__clkbuf_1 _11622_ (.A(_05293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _11623_ (.A0(\fifo_inst.mem.rMemory[13][9] ),
    .A1(_05206_),
    .S(_05289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05294_));
 sky130_fd_sc_hd__clkbuf_1 _11624_ (.A(_05294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00258_));
 sky130_fd_sc_hd__buf_2 _11625_ (.A(_05281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05295_));
 sky130_fd_sc_hd__mux2_1 _11626_ (.A0(\fifo_inst.mem.rMemory[13][10] ),
    .A1(_05208_),
    .S(_05295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05296_));
 sky130_fd_sc_hd__clkbuf_1 _11627_ (.A(_05296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _11628_ (.A0(\fifo_inst.mem.rMemory[13][11] ),
    .A1(_05211_),
    .S(_05295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05297_));
 sky130_fd_sc_hd__clkbuf_1 _11629_ (.A(_05297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _11630_ (.A0(\fifo_inst.mem.rMemory[13][12] ),
    .A1(_05213_),
    .S(_05295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05298_));
 sky130_fd_sc_hd__clkbuf_1 _11631_ (.A(_05298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _11632_ (.A0(\fifo_inst.mem.rMemory[13][13] ),
    .A1(_05215_),
    .S(_05295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05299_));
 sky130_fd_sc_hd__clkbuf_1 _11633_ (.A(_05299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _11634_ (.A0(\fifo_inst.mem.rMemory[13][14] ),
    .A1(_05217_),
    .S(_05295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05300_));
 sky130_fd_sc_hd__clkbuf_1 _11635_ (.A(_05300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00263_));
 sky130_fd_sc_hd__buf_2 _11636_ (.A(_05281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05301_));
 sky130_fd_sc_hd__mux2_1 _11637_ (.A0(\fifo_inst.mem.rMemory[13][15] ),
    .A1(_05219_),
    .S(_05301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05302_));
 sky130_fd_sc_hd__clkbuf_1 _11638_ (.A(_05302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _11639_ (.A0(\fifo_inst.mem.rMemory[13][16] ),
    .A1(_05222_),
    .S(_05301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05303_));
 sky130_fd_sc_hd__clkbuf_1 _11640_ (.A(_05303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _11641_ (.A0(\fifo_inst.mem.rMemory[13][17] ),
    .A1(_05224_),
    .S(_05301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05304_));
 sky130_fd_sc_hd__clkbuf_1 _11642_ (.A(_05304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _11643_ (.A0(\fifo_inst.mem.rMemory[13][18] ),
    .A1(_05226_),
    .S(_05301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05305_));
 sky130_fd_sc_hd__clkbuf_1 _11644_ (.A(_05305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _11645_ (.A0(\fifo_inst.mem.rMemory[13][19] ),
    .A1(_05228_),
    .S(_05301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05306_));
 sky130_fd_sc_hd__clkbuf_1 _11646_ (.A(_05306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _11647_ (.A0(\fifo_inst.mem.rMemory[13][20] ),
    .A1(_05230_),
    .S(_05282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05307_));
 sky130_fd_sc_hd__clkbuf_1 _11648_ (.A(_05307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _11649_ (.A0(\fifo_inst.mem.rMemory[13][21] ),
    .A1(_05232_),
    .S(_05282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05308_));
 sky130_fd_sc_hd__clkbuf_1 _11650_ (.A(_05308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _11651_ (.A0(\fifo_inst.mem.rMemory[13][22] ),
    .A1(_05234_),
    .S(_05282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05309_));
 sky130_fd_sc_hd__clkbuf_1 _11652_ (.A(_05309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _11653_ (.A0(\fifo_inst.mem.rMemory[13][23] ),
    .A1(_05236_),
    .S(_05282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05310_));
 sky130_fd_sc_hd__clkbuf_1 _11654_ (.A(_05310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00272_));
 sky130_fd_sc_hd__or3_4 _11655_ (.A(_05278_),
    .B(_05065_),
    .C(_05067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05311_));
 sky130_fd_sc_hd__nor2_8 _11656_ (.A(_05184_),
    .B(_05311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05312_));
 sky130_fd_sc_hd__buf_2 _11657_ (.A(_05312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05313_));
 sky130_fd_sc_hd__buf_2 _11658_ (.A(_05313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05314_));
 sky130_fd_sc_hd__mux2_1 _11659_ (.A0(\fifo_inst.mem.rMemory[12][0] ),
    .A1(_05183_),
    .S(_05314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05315_));
 sky130_fd_sc_hd__clkbuf_1 _11660_ (.A(_05315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _11661_ (.A0(\fifo_inst.mem.rMemory[12][1] ),
    .A1(_05189_),
    .S(_05314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05316_));
 sky130_fd_sc_hd__clkbuf_1 _11662_ (.A(_05316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _11663_ (.A0(\fifo_inst.mem.rMemory[12][2] ),
    .A1(_05191_),
    .S(_05314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05317_));
 sky130_fd_sc_hd__clkbuf_1 _11664_ (.A(_05317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _11665_ (.A0(\fifo_inst.mem.rMemory[12][3] ),
    .A1(_05193_),
    .S(_05314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05318_));
 sky130_fd_sc_hd__clkbuf_1 _11666_ (.A(_05318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _11667_ (.A0(\fifo_inst.mem.rMemory[12][4] ),
    .A1(_05195_),
    .S(_05314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05319_));
 sky130_fd_sc_hd__clkbuf_1 _11668_ (.A(_05319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00277_));
 sky130_fd_sc_hd__buf_2 _11669_ (.A(_05312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05320_));
 sky130_fd_sc_hd__mux2_1 _11670_ (.A0(\fifo_inst.mem.rMemory[12][5] ),
    .A1(_05197_),
    .S(_05320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05321_));
 sky130_fd_sc_hd__clkbuf_1 _11671_ (.A(_05321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _11672_ (.A0(\fifo_inst.mem.rMemory[12][6] ),
    .A1(_05200_),
    .S(_05320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05322_));
 sky130_fd_sc_hd__clkbuf_1 _11673_ (.A(_05322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _11674_ (.A0(\fifo_inst.mem.rMemory[12][7] ),
    .A1(_05202_),
    .S(_05320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05323_));
 sky130_fd_sc_hd__clkbuf_1 _11675_ (.A(_05323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _11676_ (.A0(\fifo_inst.mem.rMemory[12][8] ),
    .A1(_05204_),
    .S(_05320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05324_));
 sky130_fd_sc_hd__clkbuf_1 _11677_ (.A(_05324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _11678_ (.A0(\fifo_inst.mem.rMemory[12][9] ),
    .A1(_05206_),
    .S(_05320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05325_));
 sky130_fd_sc_hd__clkbuf_1 _11679_ (.A(_05325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00282_));
 sky130_fd_sc_hd__buf_2 _11680_ (.A(_05312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05326_));
 sky130_fd_sc_hd__mux2_1 _11681_ (.A0(\fifo_inst.mem.rMemory[12][10] ),
    .A1(_05208_),
    .S(_05326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05327_));
 sky130_fd_sc_hd__clkbuf_1 _11682_ (.A(_05327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _11683_ (.A0(\fifo_inst.mem.rMemory[12][11] ),
    .A1(_05211_),
    .S(_05326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05328_));
 sky130_fd_sc_hd__clkbuf_1 _11684_ (.A(_05328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _11685_ (.A0(\fifo_inst.mem.rMemory[12][12] ),
    .A1(_05213_),
    .S(_05326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05329_));
 sky130_fd_sc_hd__clkbuf_1 _11686_ (.A(_05329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _11687_ (.A0(\fifo_inst.mem.rMemory[12][13] ),
    .A1(_05215_),
    .S(_05326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05330_));
 sky130_fd_sc_hd__clkbuf_1 _11688_ (.A(_05330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _11689_ (.A0(\fifo_inst.mem.rMemory[12][14] ),
    .A1(_05217_),
    .S(_05326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05331_));
 sky130_fd_sc_hd__clkbuf_1 _11690_ (.A(_05331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00287_));
 sky130_fd_sc_hd__buf_2 _11691_ (.A(_05312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05332_));
 sky130_fd_sc_hd__mux2_1 _11692_ (.A0(\fifo_inst.mem.rMemory[12][15] ),
    .A1(_05219_),
    .S(_05332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05333_));
 sky130_fd_sc_hd__clkbuf_1 _11693_ (.A(_05333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _11694_ (.A0(\fifo_inst.mem.rMemory[12][16] ),
    .A1(_05222_),
    .S(_05332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05334_));
 sky130_fd_sc_hd__clkbuf_1 _11695_ (.A(_05334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00289_));
 sky130_fd_sc_hd__mux2_1 _11696_ (.A0(\fifo_inst.mem.rMemory[12][17] ),
    .A1(_05224_),
    .S(_05332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05335_));
 sky130_fd_sc_hd__clkbuf_1 _11697_ (.A(_05335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00290_));
 sky130_fd_sc_hd__mux2_1 _11698_ (.A0(\fifo_inst.mem.rMemory[12][18] ),
    .A1(_05226_),
    .S(_05332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05336_));
 sky130_fd_sc_hd__clkbuf_1 _11699_ (.A(_05336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00291_));
 sky130_fd_sc_hd__mux2_1 _11700_ (.A0(\fifo_inst.mem.rMemory[12][19] ),
    .A1(_05228_),
    .S(_05332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05337_));
 sky130_fd_sc_hd__clkbuf_1 _11701_ (.A(_05337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00292_));
 sky130_fd_sc_hd__mux2_1 _11702_ (.A0(\fifo_inst.mem.rMemory[12][20] ),
    .A1(_05230_),
    .S(_05313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05338_));
 sky130_fd_sc_hd__clkbuf_1 _11703_ (.A(_05338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _11704_ (.A0(\fifo_inst.mem.rMemory[12][21] ),
    .A1(_05232_),
    .S(_05313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05339_));
 sky130_fd_sc_hd__clkbuf_1 _11705_ (.A(_05339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _11706_ (.A0(\fifo_inst.mem.rMemory[12][22] ),
    .A1(_05234_),
    .S(_05313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05340_));
 sky130_fd_sc_hd__clkbuf_1 _11707_ (.A(_05340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _11708_ (.A0(\fifo_inst.mem.rMemory[12][23] ),
    .A1(_05236_),
    .S(_05313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05341_));
 sky130_fd_sc_hd__clkbuf_1 _11709_ (.A(_05341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00296_));
 sky130_fd_sc_hd__clkbuf_2 _11710_ (.A(_05070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05342_));
 sky130_fd_sc_hd__o31a_1 _11711_ (.A1(\shift_register[10] ),
    .A2(\shift_register[9] ),
    .A3(\shift_register[11] ),
    .B1(_05066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05343_));
 sky130_fd_sc_hd__and3_2 _11712_ (.A(\fifo_inst.mem.WR1_ADDR[1] ),
    .B(_05065_),
    .C(_05343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05344_));
 sky130_fd_sc_hd__clkbuf_2 _11713_ (.A(_05069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05345_));
 sky130_fd_sc_hd__nand3b_4 _11714_ (.A_N(_05342_),
    .B(_05344_),
    .C(_05345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05346_));
 sky130_fd_sc_hd__buf_2 _11715_ (.A(_05346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05347_));
 sky130_fd_sc_hd__buf_2 _11716_ (.A(_05347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05348_));
 sky130_fd_sc_hd__mux2_1 _11717_ (.A0(_05064_),
    .A1(\fifo_inst.mem.rMemory[11][0] ),
    .S(_05348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05349_));
 sky130_fd_sc_hd__clkbuf_1 _11718_ (.A(_05349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_1 _11719_ (.A0(_05076_),
    .A1(\fifo_inst.mem.rMemory[11][1] ),
    .S(_05348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05350_));
 sky130_fd_sc_hd__clkbuf_1 _11720_ (.A(_05350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00298_));
 sky130_fd_sc_hd__mux2_1 _11721_ (.A0(_05078_),
    .A1(\fifo_inst.mem.rMemory[11][2] ),
    .S(_05348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05351_));
 sky130_fd_sc_hd__clkbuf_1 _11722_ (.A(_05351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00299_));
 sky130_fd_sc_hd__mux2_1 _11723_ (.A0(_05080_),
    .A1(\fifo_inst.mem.rMemory[11][3] ),
    .S(_05348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05352_));
 sky130_fd_sc_hd__clkbuf_1 _11724_ (.A(_05352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _11725_ (.A0(_05082_),
    .A1(\fifo_inst.mem.rMemory[11][4] ),
    .S(_05348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05353_));
 sky130_fd_sc_hd__clkbuf_1 _11726_ (.A(_05353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00301_));
 sky130_fd_sc_hd__clkbuf_2 _11727_ (.A(_05346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05354_));
 sky130_fd_sc_hd__mux2_1 _11728_ (.A0(_05084_),
    .A1(\fifo_inst.mem.rMemory[11][5] ),
    .S(_05354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05355_));
 sky130_fd_sc_hd__clkbuf_1 _11729_ (.A(_05355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00302_));
 sky130_fd_sc_hd__mux2_1 _11730_ (.A0(_05087_),
    .A1(\fifo_inst.mem.rMemory[11][6] ),
    .S(_05354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05356_));
 sky130_fd_sc_hd__clkbuf_1 _11731_ (.A(_05356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00303_));
 sky130_fd_sc_hd__mux2_1 _11732_ (.A0(_05089_),
    .A1(\fifo_inst.mem.rMemory[11][7] ),
    .S(_05354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05357_));
 sky130_fd_sc_hd__clkbuf_1 _11733_ (.A(_05357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00304_));
 sky130_fd_sc_hd__mux2_1 _11734_ (.A0(_05091_),
    .A1(\fifo_inst.mem.rMemory[11][8] ),
    .S(_05354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05358_));
 sky130_fd_sc_hd__clkbuf_1 _11735_ (.A(_05358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00305_));
 sky130_fd_sc_hd__mux2_1 _11736_ (.A0(_05093_),
    .A1(\fifo_inst.mem.rMemory[11][9] ),
    .S(_05354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05359_));
 sky130_fd_sc_hd__clkbuf_1 _11737_ (.A(_05359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00306_));
 sky130_fd_sc_hd__buf_2 _11738_ (.A(_05346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05360_));
 sky130_fd_sc_hd__mux2_1 _11739_ (.A0(_05095_),
    .A1(\fifo_inst.mem.rMemory[11][10] ),
    .S(_05360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05361_));
 sky130_fd_sc_hd__clkbuf_1 _11740_ (.A(_05361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00307_));
 sky130_fd_sc_hd__mux2_1 _11741_ (.A0(_05098_),
    .A1(\fifo_inst.mem.rMemory[11][11] ),
    .S(_05360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05362_));
 sky130_fd_sc_hd__clkbuf_1 _11742_ (.A(_05362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_1 _11743_ (.A0(_05100_),
    .A1(\fifo_inst.mem.rMemory[11][12] ),
    .S(_05360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05363_));
 sky130_fd_sc_hd__clkbuf_1 _11744_ (.A(_05363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00309_));
 sky130_fd_sc_hd__mux2_1 _11745_ (.A0(_05102_),
    .A1(\fifo_inst.mem.rMemory[11][13] ),
    .S(_05360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05364_));
 sky130_fd_sc_hd__clkbuf_1 _11746_ (.A(_05364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00310_));
 sky130_fd_sc_hd__mux2_1 _11747_ (.A0(_05104_),
    .A1(\fifo_inst.mem.rMemory[11][14] ),
    .S(_05360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05365_));
 sky130_fd_sc_hd__clkbuf_1 _11748_ (.A(_05365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00311_));
 sky130_fd_sc_hd__clkbuf_4 _11749_ (.A(_05346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05366_));
 sky130_fd_sc_hd__mux2_1 _11750_ (.A0(_05106_),
    .A1(\fifo_inst.mem.rMemory[11][15] ),
    .S(_05366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05367_));
 sky130_fd_sc_hd__clkbuf_1 _11751_ (.A(_05367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_1 _11752_ (.A0(_05113_),
    .A1(\fifo_inst.mem.rMemory[11][16] ),
    .S(_05366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05368_));
 sky130_fd_sc_hd__clkbuf_1 _11753_ (.A(_05368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _11754_ (.A0(_05118_),
    .A1(\fifo_inst.mem.rMemory[11][17] ),
    .S(_05366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05369_));
 sky130_fd_sc_hd__clkbuf_1 _11755_ (.A(_05369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _11756_ (.A0(_05122_),
    .A1(\fifo_inst.mem.rMemory[11][18] ),
    .S(_05366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05370_));
 sky130_fd_sc_hd__clkbuf_1 _11757_ (.A(_05370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_1 _11758_ (.A0(_05127_),
    .A1(\fifo_inst.mem.rMemory[11][19] ),
    .S(_05366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05371_));
 sky130_fd_sc_hd__clkbuf_1 _11759_ (.A(_05371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _11760_ (.A0(_05131_),
    .A1(\fifo_inst.mem.rMemory[11][20] ),
    .S(_05347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05372_));
 sky130_fd_sc_hd__clkbuf_1 _11761_ (.A(_05372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _11762_ (.A0(_05136_),
    .A1(\fifo_inst.mem.rMemory[11][21] ),
    .S(_05347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05373_));
 sky130_fd_sc_hd__clkbuf_1 _11763_ (.A(_05373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _11764_ (.A0(_05140_),
    .A1(\fifo_inst.mem.rMemory[11][22] ),
    .S(_05347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05374_));
 sky130_fd_sc_hd__clkbuf_1 _11765_ (.A(_05374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_1 _11766_ (.A0(_05144_),
    .A1(\fifo_inst.mem.rMemory[11][23] ),
    .S(_05347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05375_));
 sky130_fd_sc_hd__clkbuf_1 _11767_ (.A(_05375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00320_));
 sky130_fd_sc_hd__and2_1 _11768_ (.A(\sa_inst._12_[1] ),
    .B(_00802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05376_));
 sky130_fd_sc_hd__clkbuf_1 _11769_ (.A(_05376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00321_));
 sky130_fd_sc_hd__and2_1 _11770_ (.A(\sa_inst._12_[2] ),
    .B(_00802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05377_));
 sky130_fd_sc_hd__clkbuf_1 _11771_ (.A(_05377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00322_));
 sky130_fd_sc_hd__and2_1 _11772_ (.A(\sa_inst._12_[3] ),
    .B(_00802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05378_));
 sky130_fd_sc_hd__clkbuf_1 _11773_ (.A(_05378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00323_));
 sky130_fd_sc_hd__clkbuf_2 _11774_ (.A(_00801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05379_));
 sky130_fd_sc_hd__clkbuf_1 _11775_ (.A(_05379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05380_));
 sky130_fd_sc_hd__and2_1 _11776_ (.A(\sa_inst._12_[4] ),
    .B(_05380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05381_));
 sky130_fd_sc_hd__clkbuf_1 _11777_ (.A(_05381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00324_));
 sky130_fd_sc_hd__and2_1 _11778_ (.A(\sa_inst._12_[5] ),
    .B(_05380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05382_));
 sky130_fd_sc_hd__clkbuf_1 _11779_ (.A(_05382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00325_));
 sky130_fd_sc_hd__and2_1 _11780_ (.A(\sa_inst._12_[6] ),
    .B(_05380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05383_));
 sky130_fd_sc_hd__clkbuf_1 _11781_ (.A(_05383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00326_));
 sky130_fd_sc_hd__and2_1 _11782_ (.A(\sa_inst._12_[7] ),
    .B(_05380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05384_));
 sky130_fd_sc_hd__clkbuf_1 _11783_ (.A(_05384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00327_));
 sky130_fd_sc_hd__and2_1 _11784_ (.A(\sa_inst._12_[8] ),
    .B(_05380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05385_));
 sky130_fd_sc_hd__clkbuf_1 _11785_ (.A(_05385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00328_));
 sky130_fd_sc_hd__clkbuf_1 _11786_ (.A(_05379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05386_));
 sky130_fd_sc_hd__and2_1 _11787_ (.A(\sa_inst._12_[9] ),
    .B(_05386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05387_));
 sky130_fd_sc_hd__clkbuf_1 _11788_ (.A(_05387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00329_));
 sky130_fd_sc_hd__and2_1 _11789_ (.A(\sa_inst._12_[10] ),
    .B(_05386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05388_));
 sky130_fd_sc_hd__clkbuf_1 _11790_ (.A(_05388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00330_));
 sky130_fd_sc_hd__and2_1 _11791_ (.A(\sa_inst._12_[11] ),
    .B(_05386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05389_));
 sky130_fd_sc_hd__clkbuf_1 _11792_ (.A(_05389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00331_));
 sky130_fd_sc_hd__and2_1 _11793_ (.A(\sa_inst._12_[12] ),
    .B(_05386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05390_));
 sky130_fd_sc_hd__clkbuf_1 _11794_ (.A(_05390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00332_));
 sky130_fd_sc_hd__and2_1 _11795_ (.A(\sa_inst._12_[13] ),
    .B(_05386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05391_));
 sky130_fd_sc_hd__clkbuf_1 _11796_ (.A(_05391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00333_));
 sky130_fd_sc_hd__clkbuf_1 _11797_ (.A(_00801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05392_));
 sky130_fd_sc_hd__and2_1 _11798_ (.A(\sa_inst._12_[14] ),
    .B(_05392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05393_));
 sky130_fd_sc_hd__clkbuf_1 _11799_ (.A(_05393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00334_));
 sky130_fd_sc_hd__and2_1 _11800_ (.A(\sa_inst._12_[15] ),
    .B(_05392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05394_));
 sky130_fd_sc_hd__clkbuf_1 _11801_ (.A(_05394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00335_));
 sky130_fd_sc_hd__and2_1 _11802_ (.A(\sa_inst._12_[16] ),
    .B(_05392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05395_));
 sky130_fd_sc_hd__clkbuf_1 _11803_ (.A(_05395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00336_));
 sky130_fd_sc_hd__and2_1 _11804_ (.A(\sa_inst._12_[17] ),
    .B(_05392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05396_));
 sky130_fd_sc_hd__clkbuf_1 _11805_ (.A(_05396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00337_));
 sky130_fd_sc_hd__and2_1 _11806_ (.A(\sa_inst._12_[18] ),
    .B(_05392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05397_));
 sky130_fd_sc_hd__clkbuf_1 _11807_ (.A(_05397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00338_));
 sky130_fd_sc_hd__clkbuf_1 _11808_ (.A(_00801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05398_));
 sky130_fd_sc_hd__and2_1 _11809_ (.A(\sa_inst._12_[19] ),
    .B(_05398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05399_));
 sky130_fd_sc_hd__clkbuf_1 _11810_ (.A(_05399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00339_));
 sky130_fd_sc_hd__and2_1 _11811_ (.A(\sa_inst._12_[20] ),
    .B(_05398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05400_));
 sky130_fd_sc_hd__clkbuf_1 _11812_ (.A(_05400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00340_));
 sky130_fd_sc_hd__and2_1 _11813_ (.A(\sa_inst._12_[21] ),
    .B(_05398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05401_));
 sky130_fd_sc_hd__clkbuf_1 _11814_ (.A(_05401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00341_));
 sky130_fd_sc_hd__and2_1 _11815_ (.A(\sa_inst._12_[22] ),
    .B(_05398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05402_));
 sky130_fd_sc_hd__clkbuf_1 _11816_ (.A(_05402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00342_));
 sky130_fd_sc_hd__and2_1 _11817_ (.A(\sa_inst._12_[23] ),
    .B(_05398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05403_));
 sky130_fd_sc_hd__clkbuf_1 _11818_ (.A(_05403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00343_));
 sky130_fd_sc_hd__clkbuf_1 _11819_ (.A(_00801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05404_));
 sky130_fd_sc_hd__and2_1 _11820_ (.A(\sa_inst._12_[24] ),
    .B(_05404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05405_));
 sky130_fd_sc_hd__clkbuf_1 _11821_ (.A(_05405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00344_));
 sky130_fd_sc_hd__and2_1 _11822_ (.A(\sa_inst._12_[25] ),
    .B(_05404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05406_));
 sky130_fd_sc_hd__clkbuf_1 _11823_ (.A(_05406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00345_));
 sky130_fd_sc_hd__and2_1 _11824_ (.A(\sa_inst._12_[26] ),
    .B(_05404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05407_));
 sky130_fd_sc_hd__clkbuf_1 _11825_ (.A(_05407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00346_));
 sky130_fd_sc_hd__and2_1 _11826_ (.A(\sa_inst._12_[27] ),
    .B(_05404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05408_));
 sky130_fd_sc_hd__clkbuf_1 _11827_ (.A(_05408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00347_));
 sky130_fd_sc_hd__and2_1 _11828_ (.A(\sa_inst._12_[28] ),
    .B(_05404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05409_));
 sky130_fd_sc_hd__clkbuf_1 _11829_ (.A(_05409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00348_));
 sky130_fd_sc_hd__and2_1 _11830_ (.A(\sa_inst._12_[29] ),
    .B(_05379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05410_));
 sky130_fd_sc_hd__clkbuf_1 _11831_ (.A(_05410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00349_));
 sky130_fd_sc_hd__and2_1 _11832_ (.A(\sa_inst._12_[30] ),
    .B(_05379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05411_));
 sky130_fd_sc_hd__clkbuf_1 _11833_ (.A(_05411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00350_));
 sky130_fd_sc_hd__and2_1 _11834_ (.A(\sa_inst._12_[31] ),
    .B(_05379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05412_));
 sky130_fd_sc_hd__clkbuf_1 _11835_ (.A(_05412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00351_));
 sky130_fd_sc_hd__and2_1 _11836_ (.A(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._03_ ),
    .B(_00908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05413_));
 sky130_fd_sc_hd__clkbuf_1 _11837_ (.A(_05413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00352_));
 sky130_fd_sc_hd__or4_1 _11838_ (.A(\sa_inst.cols_l2a:2.l2a_i._29_[0] ),
    .B(\sa_inst.cols_l2a:2.l2a_i._29_[1] ),
    .C(\sa_inst.cols_l2a:2.l2a_i._29_[3] ),
    .D(\sa_inst.cols_l2a:2.l2a_i._29_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05414_));
 sky130_fd_sc_hd__or4b_1 _11839_ (.A(\sa_inst.cols_l2a:2.l2a_i._29_[2] ),
    .B(\sa_inst.cols_l2a:2.l2a_i._29_[4] ),
    .C(_05414_),
    .D_N(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._55_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05415_));
 sky130_fd_sc_hd__inv_2 _11840_ (.A(_05415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00353_));
 sky130_fd_sc_hd__or2b_4 _11841_ (.A(_05070_),
    .B_N(_05069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05416_));
 sky130_fd_sc_hd__nor2_8 _11842_ (.A(_05068_),
    .B(_05416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05417_));
 sky130_fd_sc_hd__buf_2 _11843_ (.A(_05417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05418_));
 sky130_fd_sc_hd__buf_2 _11844_ (.A(_05418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05419_));
 sky130_fd_sc_hd__mux2_1 _11845_ (.A0(\fifo_inst.mem.rMemory[10][0] ),
    .A1(_05183_),
    .S(_05419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05420_));
 sky130_fd_sc_hd__clkbuf_1 _11846_ (.A(_05420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _11847_ (.A0(\fifo_inst.mem.rMemory[10][1] ),
    .A1(_05189_),
    .S(_05419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05421_));
 sky130_fd_sc_hd__clkbuf_1 _11848_ (.A(_05421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _11849_ (.A0(\fifo_inst.mem.rMemory[10][2] ),
    .A1(_05191_),
    .S(_05419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05422_));
 sky130_fd_sc_hd__clkbuf_1 _11850_ (.A(_05422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _11851_ (.A0(\fifo_inst.mem.rMemory[10][3] ),
    .A1(_05193_),
    .S(_05419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05423_));
 sky130_fd_sc_hd__clkbuf_1 _11852_ (.A(_05423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _11853_ (.A0(\fifo_inst.mem.rMemory[10][4] ),
    .A1(_05195_),
    .S(_05419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05424_));
 sky130_fd_sc_hd__clkbuf_1 _11854_ (.A(_05424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00358_));
 sky130_fd_sc_hd__clkbuf_2 _11855_ (.A(_05417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05425_));
 sky130_fd_sc_hd__mux2_1 _11856_ (.A0(\fifo_inst.mem.rMemory[10][5] ),
    .A1(_05197_),
    .S(_05425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05426_));
 sky130_fd_sc_hd__clkbuf_1 _11857_ (.A(_05426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _11858_ (.A0(\fifo_inst.mem.rMemory[10][6] ),
    .A1(_05200_),
    .S(_05425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05427_));
 sky130_fd_sc_hd__clkbuf_1 _11859_ (.A(_05427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _11860_ (.A0(\fifo_inst.mem.rMemory[10][7] ),
    .A1(_05202_),
    .S(_05425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05428_));
 sky130_fd_sc_hd__clkbuf_1 _11861_ (.A(_05428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _11862_ (.A0(\fifo_inst.mem.rMemory[10][8] ),
    .A1(_05204_),
    .S(_05425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05429_));
 sky130_fd_sc_hd__clkbuf_1 _11863_ (.A(_05429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _11864_ (.A0(\fifo_inst.mem.rMemory[10][9] ),
    .A1(_05206_),
    .S(_05425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05430_));
 sky130_fd_sc_hd__clkbuf_1 _11865_ (.A(_05430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00363_));
 sky130_fd_sc_hd__clkbuf_2 _11866_ (.A(_05417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05431_));
 sky130_fd_sc_hd__mux2_1 _11867_ (.A0(\fifo_inst.mem.rMemory[10][10] ),
    .A1(_05208_),
    .S(_05431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05432_));
 sky130_fd_sc_hd__clkbuf_1 _11868_ (.A(_05432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _11869_ (.A0(\fifo_inst.mem.rMemory[10][11] ),
    .A1(_05211_),
    .S(_05431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05433_));
 sky130_fd_sc_hd__clkbuf_1 _11870_ (.A(_05433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _11871_ (.A0(\fifo_inst.mem.rMemory[10][12] ),
    .A1(_05213_),
    .S(_05431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05434_));
 sky130_fd_sc_hd__clkbuf_1 _11872_ (.A(_05434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_1 _11873_ (.A0(\fifo_inst.mem.rMemory[10][13] ),
    .A1(_05215_),
    .S(_05431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05435_));
 sky130_fd_sc_hd__clkbuf_1 _11874_ (.A(_05435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _11875_ (.A0(\fifo_inst.mem.rMemory[10][14] ),
    .A1(_05217_),
    .S(_05431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05436_));
 sky130_fd_sc_hd__clkbuf_1 _11876_ (.A(_05436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00368_));
 sky130_fd_sc_hd__buf_2 _11877_ (.A(_05417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05437_));
 sky130_fd_sc_hd__mux2_1 _11878_ (.A0(\fifo_inst.mem.rMemory[10][15] ),
    .A1(_05219_),
    .S(_05437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05438_));
 sky130_fd_sc_hd__clkbuf_1 _11879_ (.A(_05438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _11880_ (.A0(\fifo_inst.mem.rMemory[10][16] ),
    .A1(_05222_),
    .S(_05437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05439_));
 sky130_fd_sc_hd__clkbuf_1 _11881_ (.A(_05439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _11882_ (.A0(\fifo_inst.mem.rMemory[10][17] ),
    .A1(_05224_),
    .S(_05437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05440_));
 sky130_fd_sc_hd__clkbuf_1 _11883_ (.A(_05440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _11884_ (.A0(\fifo_inst.mem.rMemory[10][18] ),
    .A1(_05226_),
    .S(_05437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05441_));
 sky130_fd_sc_hd__clkbuf_1 _11885_ (.A(_05441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _11886_ (.A0(\fifo_inst.mem.rMemory[10][19] ),
    .A1(_05228_),
    .S(_05437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05442_));
 sky130_fd_sc_hd__clkbuf_1 _11887_ (.A(_05442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _11888_ (.A0(\fifo_inst.mem.rMemory[10][20] ),
    .A1(_05230_),
    .S(_05418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05443_));
 sky130_fd_sc_hd__clkbuf_1 _11889_ (.A(_05443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_1 _11890_ (.A0(\fifo_inst.mem.rMemory[10][21] ),
    .A1(_05232_),
    .S(_05418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05444_));
 sky130_fd_sc_hd__clkbuf_1 _11891_ (.A(_05444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _11892_ (.A0(\fifo_inst.mem.rMemory[10][22] ),
    .A1(_05234_),
    .S(_05418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05445_));
 sky130_fd_sc_hd__clkbuf_1 _11893_ (.A(_05445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _11894_ (.A0(\fifo_inst.mem.rMemory[10][23] ),
    .A1(_05236_),
    .S(_05418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05446_));
 sky130_fd_sc_hd__clkbuf_1 _11895_ (.A(_05446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00377_));
 sky130_fd_sc_hd__nor2_8 _11896_ (.A(_05071_),
    .B(_05311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05447_));
 sky130_fd_sc_hd__clkbuf_2 _11897_ (.A(_05447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05448_));
 sky130_fd_sc_hd__buf_2 _11898_ (.A(_05448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05449_));
 sky130_fd_sc_hd__mux2_1 _11899_ (.A0(\fifo_inst.mem.rMemory[0][0] ),
    .A1(_05183_),
    .S(_05449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05450_));
 sky130_fd_sc_hd__clkbuf_1 _11900_ (.A(_05450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _11901_ (.A0(\fifo_inst.mem.rMemory[0][1] ),
    .A1(_05189_),
    .S(_05449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05451_));
 sky130_fd_sc_hd__clkbuf_1 _11902_ (.A(_05451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _11903_ (.A0(\fifo_inst.mem.rMemory[0][2] ),
    .A1(_05191_),
    .S(_05449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05452_));
 sky130_fd_sc_hd__clkbuf_1 _11904_ (.A(_05452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _11905_ (.A0(\fifo_inst.mem.rMemory[0][3] ),
    .A1(_05193_),
    .S(_05449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05453_));
 sky130_fd_sc_hd__clkbuf_1 _11906_ (.A(_05453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_1 _11907_ (.A0(\fifo_inst.mem.rMemory[0][4] ),
    .A1(_05195_),
    .S(_05449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05454_));
 sky130_fd_sc_hd__clkbuf_1 _11908_ (.A(_05454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00382_));
 sky130_fd_sc_hd__buf_2 _11909_ (.A(_05447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05455_));
 sky130_fd_sc_hd__mux2_1 _11910_ (.A0(\fifo_inst.mem.rMemory[0][5] ),
    .A1(_05197_),
    .S(_05455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05456_));
 sky130_fd_sc_hd__clkbuf_1 _11911_ (.A(_05456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_1 _11912_ (.A0(\fifo_inst.mem.rMemory[0][6] ),
    .A1(_05200_),
    .S(_05455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05457_));
 sky130_fd_sc_hd__clkbuf_1 _11913_ (.A(_05457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_1 _11914_ (.A0(\fifo_inst.mem.rMemory[0][7] ),
    .A1(_05202_),
    .S(_05455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05458_));
 sky130_fd_sc_hd__clkbuf_1 _11915_ (.A(_05458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_1 _11916_ (.A0(\fifo_inst.mem.rMemory[0][8] ),
    .A1(_05204_),
    .S(_05455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05459_));
 sky130_fd_sc_hd__clkbuf_1 _11917_ (.A(_05459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_1 _11918_ (.A0(\fifo_inst.mem.rMemory[0][9] ),
    .A1(_05206_),
    .S(_05455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05460_));
 sky130_fd_sc_hd__clkbuf_1 _11919_ (.A(_05460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00387_));
 sky130_fd_sc_hd__buf_2 _11920_ (.A(_05447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05461_));
 sky130_fd_sc_hd__mux2_1 _11921_ (.A0(\fifo_inst.mem.rMemory[0][10] ),
    .A1(_05208_),
    .S(_05461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05462_));
 sky130_fd_sc_hd__clkbuf_1 _11922_ (.A(_05462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _11923_ (.A0(\fifo_inst.mem.rMemory[0][11] ),
    .A1(_05211_),
    .S(_05461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05463_));
 sky130_fd_sc_hd__clkbuf_1 _11924_ (.A(_05463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _11925_ (.A0(\fifo_inst.mem.rMemory[0][12] ),
    .A1(_05213_),
    .S(_05461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05464_));
 sky130_fd_sc_hd__clkbuf_1 _11926_ (.A(_05464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00390_));
 sky130_fd_sc_hd__mux2_1 _11927_ (.A0(\fifo_inst.mem.rMemory[0][13] ),
    .A1(_05215_),
    .S(_05461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05465_));
 sky130_fd_sc_hd__clkbuf_1 _11928_ (.A(_05465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_1 _11929_ (.A0(\fifo_inst.mem.rMemory[0][14] ),
    .A1(_05217_),
    .S(_05461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05466_));
 sky130_fd_sc_hd__clkbuf_1 _11930_ (.A(_05466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00392_));
 sky130_fd_sc_hd__buf_2 _11931_ (.A(_05447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05467_));
 sky130_fd_sc_hd__mux2_1 _11932_ (.A0(\fifo_inst.mem.rMemory[0][15] ),
    .A1(_05219_),
    .S(_05467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05468_));
 sky130_fd_sc_hd__clkbuf_1 _11933_ (.A(_05468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00393_));
 sky130_fd_sc_hd__mux2_1 _11934_ (.A0(\fifo_inst.mem.rMemory[0][16] ),
    .A1(_05222_),
    .S(_05467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05469_));
 sky130_fd_sc_hd__clkbuf_1 _11935_ (.A(_05469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00394_));
 sky130_fd_sc_hd__mux2_1 _11936_ (.A0(\fifo_inst.mem.rMemory[0][17] ),
    .A1(_05224_),
    .S(_05467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05470_));
 sky130_fd_sc_hd__clkbuf_1 _11937_ (.A(_05470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_1 _11938_ (.A0(\fifo_inst.mem.rMemory[0][18] ),
    .A1(_05226_),
    .S(_05467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05471_));
 sky130_fd_sc_hd__clkbuf_1 _11939_ (.A(_05471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00396_));
 sky130_fd_sc_hd__mux2_1 _11940_ (.A0(\fifo_inst.mem.rMemory[0][19] ),
    .A1(_05228_),
    .S(_05467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05472_));
 sky130_fd_sc_hd__clkbuf_1 _11941_ (.A(_05472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _11942_ (.A0(\fifo_inst.mem.rMemory[0][20] ),
    .A1(_05230_),
    .S(_05448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05473_));
 sky130_fd_sc_hd__clkbuf_1 _11943_ (.A(_05473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_1 _11944_ (.A0(\fifo_inst.mem.rMemory[0][21] ),
    .A1(_05232_),
    .S(_05448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05474_));
 sky130_fd_sc_hd__clkbuf_1 _11945_ (.A(_05474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_1 _11946_ (.A0(\fifo_inst.mem.rMemory[0][22] ),
    .A1(_05234_),
    .S(_05448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05475_));
 sky130_fd_sc_hd__clkbuf_1 _11947_ (.A(_05475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00400_));
 sky130_fd_sc_hd__mux2_1 _11948_ (.A0(\fifo_inst.mem.rMemory[0][23] ),
    .A1(_05236_),
    .S(_05448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05476_));
 sky130_fd_sc_hd__clkbuf_1 _11949_ (.A(_05476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00401_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11950_ (.A(\fifo_inst.WR_DATA[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05477_));
 sky130_fd_sc_hd__nor2_4 _11951_ (.A(_05311_),
    .B(_05416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05478_));
 sky130_fd_sc_hd__buf_2 _11952_ (.A(_05478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05479_));
 sky130_fd_sc_hd__buf_2 _11953_ (.A(_05479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05480_));
 sky130_fd_sc_hd__mux2_1 _11954_ (.A0(\fifo_inst.mem.rMemory[8][0] ),
    .A1(_05477_),
    .S(_05480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05481_));
 sky130_fd_sc_hd__clkbuf_1 _11955_ (.A(_05481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00402_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11956_ (.A(\fifo_inst.WR_DATA[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05482_));
 sky130_fd_sc_hd__mux2_1 _11957_ (.A0(\fifo_inst.mem.rMemory[8][1] ),
    .A1(_05482_),
    .S(_05480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05483_));
 sky130_fd_sc_hd__clkbuf_1 _11958_ (.A(_05483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00403_));
 sky130_fd_sc_hd__clkbuf_2 _11959_ (.A(\fifo_inst.WR_DATA[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05484_));
 sky130_fd_sc_hd__mux2_1 _11960_ (.A0(\fifo_inst.mem.rMemory[8][2] ),
    .A1(_05484_),
    .S(_05480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05485_));
 sky130_fd_sc_hd__clkbuf_1 _11961_ (.A(_05485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00404_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11962_ (.A(\fifo_inst.WR_DATA[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05486_));
 sky130_fd_sc_hd__mux2_1 _11963_ (.A0(\fifo_inst.mem.rMemory[8][3] ),
    .A1(_05486_),
    .S(_05480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05487_));
 sky130_fd_sc_hd__clkbuf_1 _11964_ (.A(_05487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00405_));
 sky130_fd_sc_hd__clkbuf_2 _11965_ (.A(\fifo_inst.WR_DATA[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05488_));
 sky130_fd_sc_hd__mux2_1 _11966_ (.A0(\fifo_inst.mem.rMemory[8][4] ),
    .A1(_05488_),
    .S(_05480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05489_));
 sky130_fd_sc_hd__clkbuf_1 _11967_ (.A(_05489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00406_));
 sky130_fd_sc_hd__clkbuf_2 _11968_ (.A(\fifo_inst.WR_DATA[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05490_));
 sky130_fd_sc_hd__clkbuf_2 _11969_ (.A(_05478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05491_));
 sky130_fd_sc_hd__mux2_1 _11970_ (.A0(\fifo_inst.mem.rMemory[8][5] ),
    .A1(_05490_),
    .S(_05491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05492_));
 sky130_fd_sc_hd__clkbuf_1 _11971_ (.A(_05492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00407_));
 sky130_fd_sc_hd__clkbuf_2 _11972_ (.A(\fifo_inst.WR_DATA[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05493_));
 sky130_fd_sc_hd__mux2_1 _11973_ (.A0(\fifo_inst.mem.rMemory[8][6] ),
    .A1(_05493_),
    .S(_05491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05494_));
 sky130_fd_sc_hd__clkbuf_1 _11974_ (.A(_05494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00408_));
 sky130_fd_sc_hd__clkbuf_2 _11975_ (.A(\fifo_inst.WR_DATA[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05495_));
 sky130_fd_sc_hd__mux2_1 _11976_ (.A0(\fifo_inst.mem.rMemory[8][7] ),
    .A1(_05495_),
    .S(_05491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05496_));
 sky130_fd_sc_hd__clkbuf_1 _11977_ (.A(_05496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00409_));
 sky130_fd_sc_hd__clkbuf_2 _11978_ (.A(\fifo_inst.WR_DATA[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05497_));
 sky130_fd_sc_hd__mux2_1 _11979_ (.A0(\fifo_inst.mem.rMemory[8][8] ),
    .A1(_05497_),
    .S(_05491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05498_));
 sky130_fd_sc_hd__clkbuf_1 _11980_ (.A(_05498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00410_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11981_ (.A(\fifo_inst.WR_DATA[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05499_));
 sky130_fd_sc_hd__mux2_1 _11982_ (.A0(\fifo_inst.mem.rMemory[8][9] ),
    .A1(_05499_),
    .S(_05491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05500_));
 sky130_fd_sc_hd__clkbuf_1 _11983_ (.A(_05500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00411_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11984_ (.A(\fifo_inst.WR_DATA[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05501_));
 sky130_fd_sc_hd__buf_2 _11985_ (.A(_05478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05502_));
 sky130_fd_sc_hd__mux2_1 _11986_ (.A0(\fifo_inst.mem.rMemory[8][10] ),
    .A1(_05501_),
    .S(_05502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05503_));
 sky130_fd_sc_hd__clkbuf_1 _11987_ (.A(_05503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00412_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11988_ (.A(\fifo_inst.WR_DATA[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05504_));
 sky130_fd_sc_hd__mux2_1 _11989_ (.A0(\fifo_inst.mem.rMemory[8][11] ),
    .A1(_05504_),
    .S(_05502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05505_));
 sky130_fd_sc_hd__clkbuf_1 _11990_ (.A(_05505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00413_));
 sky130_fd_sc_hd__clkbuf_2 _11991_ (.A(\fifo_inst.WR_DATA[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05506_));
 sky130_fd_sc_hd__mux2_1 _11992_ (.A0(\fifo_inst.mem.rMemory[8][12] ),
    .A1(_05506_),
    .S(_05502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05507_));
 sky130_fd_sc_hd__clkbuf_1 _11993_ (.A(_05507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00414_));
 sky130_fd_sc_hd__buf_2 _11994_ (.A(\fifo_inst.WR_DATA[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05508_));
 sky130_fd_sc_hd__mux2_1 _11995_ (.A0(\fifo_inst.mem.rMemory[8][13] ),
    .A1(_05508_),
    .S(_05502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05509_));
 sky130_fd_sc_hd__clkbuf_1 _11996_ (.A(_05509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00415_));
 sky130_fd_sc_hd__clkbuf_2 _11997_ (.A(\fifo_inst.WR_DATA[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05510_));
 sky130_fd_sc_hd__mux2_1 _11998_ (.A0(\fifo_inst.mem.rMemory[8][14] ),
    .A1(_05510_),
    .S(_05502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05511_));
 sky130_fd_sc_hd__clkbuf_1 _11999_ (.A(_05511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00416_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12000_ (.A(\fifo_inst.WR_DATA[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05512_));
 sky130_fd_sc_hd__clkbuf_4 _12001_ (.A(_05478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05513_));
 sky130_fd_sc_hd__mux2_1 _12002_ (.A0(\fifo_inst.mem.rMemory[8][15] ),
    .A1(_05512_),
    .S(_05513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05514_));
 sky130_fd_sc_hd__clkbuf_1 _12003_ (.A(_05514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00417_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12004_ (.A(_05112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05515_));
 sky130_fd_sc_hd__mux2_1 _12005_ (.A0(\fifo_inst.mem.rMemory[8][16] ),
    .A1(_05515_),
    .S(_05513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05516_));
 sky130_fd_sc_hd__clkbuf_1 _12006_ (.A(_05516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00418_));
 sky130_fd_sc_hd__clkbuf_2 _12007_ (.A(_05117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05517_));
 sky130_fd_sc_hd__mux2_1 _12008_ (.A0(\fifo_inst.mem.rMemory[8][17] ),
    .A1(_05517_),
    .S(_05513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05518_));
 sky130_fd_sc_hd__clkbuf_1 _12009_ (.A(_05518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00419_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12010_ (.A(_05121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05519_));
 sky130_fd_sc_hd__mux2_1 _12011_ (.A0(\fifo_inst.mem.rMemory[8][18] ),
    .A1(_05519_),
    .S(_05513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05520_));
 sky130_fd_sc_hd__clkbuf_1 _12012_ (.A(_05520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00420_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12013_ (.A(_05126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05521_));
 sky130_fd_sc_hd__mux2_1 _12014_ (.A0(\fifo_inst.mem.rMemory[8][19] ),
    .A1(_05521_),
    .S(_05513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05522_));
 sky130_fd_sc_hd__clkbuf_1 _12015_ (.A(_05522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00421_));
 sky130_fd_sc_hd__clkbuf_2 _12016_ (.A(_05130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05523_));
 sky130_fd_sc_hd__mux2_1 _12017_ (.A0(\fifo_inst.mem.rMemory[8][20] ),
    .A1(_05523_),
    .S(_05479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05524_));
 sky130_fd_sc_hd__clkbuf_1 _12018_ (.A(_05524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00422_));
 sky130_fd_sc_hd__clkbuf_2 _12019_ (.A(_05135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05525_));
 sky130_fd_sc_hd__mux2_1 _12020_ (.A0(\fifo_inst.mem.rMemory[8][21] ),
    .A1(_05525_),
    .S(_05479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05526_));
 sky130_fd_sc_hd__clkbuf_1 _12021_ (.A(_05526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00423_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12022_ (.A(_05139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05527_));
 sky130_fd_sc_hd__mux2_1 _12023_ (.A0(\fifo_inst.mem.rMemory[8][22] ),
    .A1(_05527_),
    .S(_05479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05528_));
 sky130_fd_sc_hd__clkbuf_1 _12024_ (.A(_05528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00424_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12025_ (.A(_05143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05529_));
 sky130_fd_sc_hd__mux2_1 _12026_ (.A0(\fifo_inst.mem.rMemory[8][23] ),
    .A1(_05529_),
    .S(_05479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05530_));
 sky130_fd_sc_hd__clkbuf_1 _12027_ (.A(_05530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00425_));
 sky130_fd_sc_hd__and3_1 _12028_ (.A(\sa_inst._17_[0] ),
    .B(_01032_),
    .C(_00806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05531_));
 sky130_fd_sc_hd__clkbuf_1 _12029_ (.A(_05531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00426_));
 sky130_fd_sc_hd__and3_1 _12030_ (.A(\sa_inst._17_[1] ),
    .B(_01032_),
    .C(_00806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05532_));
 sky130_fd_sc_hd__clkbuf_1 _12031_ (.A(_05532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00427_));
 sky130_fd_sc_hd__and2_1 _12032_ (.A(\sa_inst._17_[2] ),
    .B(_01032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05533_));
 sky130_fd_sc_hd__clkbuf_1 _12033_ (.A(_05533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00428_));
 sky130_fd_sc_hd__and2_1 _12034_ (.A(\sa_inst._17_[3] ),
    .B(_01032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05534_));
 sky130_fd_sc_hd__clkbuf_1 _12035_ (.A(_05534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00429_));
 sky130_fd_sc_hd__and2_1 _12036_ (.A(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._03_ ),
    .B(_00958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05535_));
 sky130_fd_sc_hd__clkbuf_1 _12037_ (.A(_05535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00430_));
 sky130_fd_sc_hd__or4_1 _12038_ (.A(\sa_inst.cols_l2a:1.l2a_i._29_[0] ),
    .B(\sa_inst.cols_l2a:1.l2a_i._29_[1] ),
    .C(\sa_inst.cols_l2a:1.l2a_i._29_[3] ),
    .D(\sa_inst.cols_l2a:1.l2a_i._29_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05536_));
 sky130_fd_sc_hd__or4b_1 _12039_ (.A(\sa_inst.cols_l2a:1.l2a_i._29_[2] ),
    .B(\sa_inst.cols_l2a:1.l2a_i._29_[4] ),
    .C(_05536_),
    .D_N(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._55_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05537_));
 sky130_fd_sc_hd__inv_2 _12040_ (.A(_05537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00431_));
 sky130_fd_sc_hd__nand3b_4 _12041_ (.A_N(_05345_),
    .B(_05342_),
    .C(_05344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05538_));
 sky130_fd_sc_hd__buf_2 _12042_ (.A(_05538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05539_));
 sky130_fd_sc_hd__buf_2 _12043_ (.A(_05539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05540_));
 sky130_fd_sc_hd__mux2_1 _12044_ (.A0(_05064_),
    .A1(\fifo_inst.mem.rMemory[7][0] ),
    .S(_05540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05541_));
 sky130_fd_sc_hd__clkbuf_1 _12045_ (.A(_05541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_1 _12046_ (.A0(_05076_),
    .A1(\fifo_inst.mem.rMemory[7][1] ),
    .S(_05540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05542_));
 sky130_fd_sc_hd__clkbuf_1 _12047_ (.A(_05542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_1 _12048_ (.A0(_05078_),
    .A1(\fifo_inst.mem.rMemory[7][2] ),
    .S(_05540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05543_));
 sky130_fd_sc_hd__clkbuf_1 _12049_ (.A(_05543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_1 _12050_ (.A0(_05080_),
    .A1(\fifo_inst.mem.rMemory[7][3] ),
    .S(_05540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05544_));
 sky130_fd_sc_hd__clkbuf_1 _12051_ (.A(_05544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _12052_ (.A0(_05082_),
    .A1(\fifo_inst.mem.rMemory[7][4] ),
    .S(_05540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05545_));
 sky130_fd_sc_hd__clkbuf_1 _12053_ (.A(_05545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00436_));
 sky130_fd_sc_hd__clkbuf_2 _12054_ (.A(_05538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05546_));
 sky130_fd_sc_hd__mux2_1 _12055_ (.A0(_05084_),
    .A1(\fifo_inst.mem.rMemory[7][5] ),
    .S(_05546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05547_));
 sky130_fd_sc_hd__clkbuf_1 _12056_ (.A(_05547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _12057_ (.A0(_05087_),
    .A1(\fifo_inst.mem.rMemory[7][6] ),
    .S(_05546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05548_));
 sky130_fd_sc_hd__clkbuf_1 _12058_ (.A(_05548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _12059_ (.A0(_05089_),
    .A1(\fifo_inst.mem.rMemory[7][7] ),
    .S(_05546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05549_));
 sky130_fd_sc_hd__clkbuf_1 _12060_ (.A(_05549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _12061_ (.A0(_05091_),
    .A1(\fifo_inst.mem.rMemory[7][8] ),
    .S(_05546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05550_));
 sky130_fd_sc_hd__clkbuf_1 _12062_ (.A(_05550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _12063_ (.A0(_05093_),
    .A1(\fifo_inst.mem.rMemory[7][9] ),
    .S(_05546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05551_));
 sky130_fd_sc_hd__clkbuf_1 _12064_ (.A(_05551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00441_));
 sky130_fd_sc_hd__buf_2 _12065_ (.A(_05538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05552_));
 sky130_fd_sc_hd__mux2_1 _12066_ (.A0(_05095_),
    .A1(\fifo_inst.mem.rMemory[7][10] ),
    .S(_05552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05553_));
 sky130_fd_sc_hd__clkbuf_1 _12067_ (.A(_05553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _12068_ (.A0(_05098_),
    .A1(\fifo_inst.mem.rMemory[7][11] ),
    .S(_05552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05554_));
 sky130_fd_sc_hd__clkbuf_1 _12069_ (.A(_05554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _12070_ (.A0(_05100_),
    .A1(\fifo_inst.mem.rMemory[7][12] ),
    .S(_05552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05555_));
 sky130_fd_sc_hd__clkbuf_1 _12071_ (.A(_05555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _12072_ (.A0(_05102_),
    .A1(\fifo_inst.mem.rMemory[7][13] ),
    .S(_05552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05556_));
 sky130_fd_sc_hd__clkbuf_1 _12073_ (.A(_05556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _12074_ (.A0(_05104_),
    .A1(\fifo_inst.mem.rMemory[7][14] ),
    .S(_05552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05557_));
 sky130_fd_sc_hd__clkbuf_1 _12075_ (.A(_05557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00446_));
 sky130_fd_sc_hd__buf_2 _12076_ (.A(_05538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05558_));
 sky130_fd_sc_hd__mux2_1 _12077_ (.A0(_05106_),
    .A1(\fifo_inst.mem.rMemory[7][15] ),
    .S(_05558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05559_));
 sky130_fd_sc_hd__clkbuf_1 _12078_ (.A(_05559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _12079_ (.A0(_05113_),
    .A1(\fifo_inst.mem.rMemory[7][16] ),
    .S(_05558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05560_));
 sky130_fd_sc_hd__clkbuf_1 _12080_ (.A(_05560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _12081_ (.A0(_05118_),
    .A1(\fifo_inst.mem.rMemory[7][17] ),
    .S(_05558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05561_));
 sky130_fd_sc_hd__clkbuf_1 _12082_ (.A(_05561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _12083_ (.A0(_05122_),
    .A1(\fifo_inst.mem.rMemory[7][18] ),
    .S(_05558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05562_));
 sky130_fd_sc_hd__clkbuf_1 _12084_ (.A(_05562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _12085_ (.A0(_05127_),
    .A1(\fifo_inst.mem.rMemory[7][19] ),
    .S(_05558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05563_));
 sky130_fd_sc_hd__clkbuf_1 _12086_ (.A(_05563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _12087_ (.A0(_05131_),
    .A1(\fifo_inst.mem.rMemory[7][20] ),
    .S(_05539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05564_));
 sky130_fd_sc_hd__clkbuf_1 _12088_ (.A(_05564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _12089_ (.A0(_05136_),
    .A1(\fifo_inst.mem.rMemory[7][21] ),
    .S(_05539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05565_));
 sky130_fd_sc_hd__clkbuf_1 _12090_ (.A(_05565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _12091_ (.A0(_05140_),
    .A1(\fifo_inst.mem.rMemory[7][22] ),
    .S(_05539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05566_));
 sky130_fd_sc_hd__clkbuf_1 _12092_ (.A(_05566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _12093_ (.A0(_05144_),
    .A1(\fifo_inst.mem.rMemory[7][23] ),
    .S(_05539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05567_));
 sky130_fd_sc_hd__clkbuf_1 _12094_ (.A(_05567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00455_));
 sky130_fd_sc_hd__nor2_4 _12095_ (.A(_05280_),
    .B(_05416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05568_));
 sky130_fd_sc_hd__buf_2 _12096_ (.A(_05568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05569_));
 sky130_fd_sc_hd__buf_2 _12097_ (.A(_05569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05570_));
 sky130_fd_sc_hd__mux2_1 _12098_ (.A0(\fifo_inst.mem.rMemory[9][0] ),
    .A1(_05477_),
    .S(_05570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05571_));
 sky130_fd_sc_hd__clkbuf_1 _12099_ (.A(_05571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _12100_ (.A0(\fifo_inst.mem.rMemory[9][1] ),
    .A1(_05482_),
    .S(_05570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05572_));
 sky130_fd_sc_hd__clkbuf_1 _12101_ (.A(_05572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _12102_ (.A0(\fifo_inst.mem.rMemory[9][2] ),
    .A1(_05484_),
    .S(_05570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05573_));
 sky130_fd_sc_hd__clkbuf_1 _12103_ (.A(_05573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _12104_ (.A0(\fifo_inst.mem.rMemory[9][3] ),
    .A1(_05486_),
    .S(_05570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05574_));
 sky130_fd_sc_hd__clkbuf_1 _12105_ (.A(_05574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _12106_ (.A0(\fifo_inst.mem.rMemory[9][4] ),
    .A1(_05488_),
    .S(_05570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05575_));
 sky130_fd_sc_hd__clkbuf_1 _12107_ (.A(_05575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00460_));
 sky130_fd_sc_hd__clkbuf_2 _12108_ (.A(_05568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05576_));
 sky130_fd_sc_hd__mux2_1 _12109_ (.A0(\fifo_inst.mem.rMemory[9][5] ),
    .A1(_05490_),
    .S(_05576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05577_));
 sky130_fd_sc_hd__clkbuf_1 _12110_ (.A(_05577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _12111_ (.A0(\fifo_inst.mem.rMemory[9][6] ),
    .A1(_05493_),
    .S(_05576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05578_));
 sky130_fd_sc_hd__clkbuf_1 _12112_ (.A(_05578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _12113_ (.A0(\fifo_inst.mem.rMemory[9][7] ),
    .A1(_05495_),
    .S(_05576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05579_));
 sky130_fd_sc_hd__clkbuf_1 _12114_ (.A(_05579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _12115_ (.A0(\fifo_inst.mem.rMemory[9][8] ),
    .A1(_05497_),
    .S(_05576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05580_));
 sky130_fd_sc_hd__clkbuf_1 _12116_ (.A(_05580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _12117_ (.A0(\fifo_inst.mem.rMemory[9][9] ),
    .A1(_05499_),
    .S(_05576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05581_));
 sky130_fd_sc_hd__clkbuf_1 _12118_ (.A(_05581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00465_));
 sky130_fd_sc_hd__buf_2 _12119_ (.A(_05568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05582_));
 sky130_fd_sc_hd__mux2_1 _12120_ (.A0(\fifo_inst.mem.rMemory[9][10] ),
    .A1(_05501_),
    .S(_05582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05583_));
 sky130_fd_sc_hd__clkbuf_1 _12121_ (.A(_05583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _12122_ (.A0(\fifo_inst.mem.rMemory[9][11] ),
    .A1(_05504_),
    .S(_05582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05584_));
 sky130_fd_sc_hd__clkbuf_1 _12123_ (.A(_05584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _12124_ (.A0(\fifo_inst.mem.rMemory[9][12] ),
    .A1(_05506_),
    .S(_05582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05585_));
 sky130_fd_sc_hd__clkbuf_1 _12125_ (.A(_05585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _12126_ (.A0(\fifo_inst.mem.rMemory[9][13] ),
    .A1(_05508_),
    .S(_05582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05586_));
 sky130_fd_sc_hd__clkbuf_1 _12127_ (.A(_05586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _12128_ (.A0(\fifo_inst.mem.rMemory[9][14] ),
    .A1(_05510_),
    .S(_05582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05587_));
 sky130_fd_sc_hd__clkbuf_1 _12129_ (.A(_05587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00470_));
 sky130_fd_sc_hd__clkbuf_4 _12130_ (.A(_05568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05588_));
 sky130_fd_sc_hd__mux2_1 _12131_ (.A0(\fifo_inst.mem.rMemory[9][15] ),
    .A1(_05512_),
    .S(_05588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05589_));
 sky130_fd_sc_hd__clkbuf_1 _12132_ (.A(_05589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _12133_ (.A0(\fifo_inst.mem.rMemory[9][16] ),
    .A1(_05515_),
    .S(_05588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05590_));
 sky130_fd_sc_hd__clkbuf_1 _12134_ (.A(_05590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _12135_ (.A0(\fifo_inst.mem.rMemory[9][17] ),
    .A1(_05517_),
    .S(_05588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05591_));
 sky130_fd_sc_hd__clkbuf_1 _12136_ (.A(_05591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _12137_ (.A0(\fifo_inst.mem.rMemory[9][18] ),
    .A1(_05519_),
    .S(_05588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05592_));
 sky130_fd_sc_hd__clkbuf_1 _12138_ (.A(_05592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _12139_ (.A0(\fifo_inst.mem.rMemory[9][19] ),
    .A1(_05521_),
    .S(_05588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05593_));
 sky130_fd_sc_hd__clkbuf_1 _12140_ (.A(_05593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _12141_ (.A0(\fifo_inst.mem.rMemory[9][20] ),
    .A1(_05523_),
    .S(_05569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05594_));
 sky130_fd_sc_hd__clkbuf_1 _12142_ (.A(_05594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _12143_ (.A0(\fifo_inst.mem.rMemory[9][21] ),
    .A1(_05525_),
    .S(_05569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05595_));
 sky130_fd_sc_hd__clkbuf_1 _12144_ (.A(_05595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _12145_ (.A0(\fifo_inst.mem.rMemory[9][22] ),
    .A1(_05527_),
    .S(_05569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05596_));
 sky130_fd_sc_hd__clkbuf_1 _12146_ (.A(_05596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _12147_ (.A0(\fifo_inst.mem.rMemory[9][23] ),
    .A1(_05529_),
    .S(_05569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05597_));
 sky130_fd_sc_hd__clkbuf_1 _12148_ (.A(_05597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00479_));
 sky130_fd_sc_hd__or2b_2 _12149_ (.A(_05069_),
    .B_N(_05070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05598_));
 sky130_fd_sc_hd__nor2_4 _12150_ (.A(_05068_),
    .B(_05598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05599_));
 sky130_fd_sc_hd__buf_2 _12151_ (.A(_05599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05600_));
 sky130_fd_sc_hd__buf_2 _12152_ (.A(_05600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05601_));
 sky130_fd_sc_hd__mux2_1 _12153_ (.A0(\fifo_inst.mem.rMemory[6][0] ),
    .A1(_05477_),
    .S(_05601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05602_));
 sky130_fd_sc_hd__clkbuf_1 _12154_ (.A(_05602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _12155_ (.A0(\fifo_inst.mem.rMemory[6][1] ),
    .A1(_05482_),
    .S(_05601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05603_));
 sky130_fd_sc_hd__clkbuf_1 _12156_ (.A(_05603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _12157_ (.A0(\fifo_inst.mem.rMemory[6][2] ),
    .A1(_05484_),
    .S(_05601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05604_));
 sky130_fd_sc_hd__clkbuf_1 _12158_ (.A(_05604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _12159_ (.A0(\fifo_inst.mem.rMemory[6][3] ),
    .A1(_05486_),
    .S(_05601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05605_));
 sky130_fd_sc_hd__clkbuf_1 _12160_ (.A(_05605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _12161_ (.A0(\fifo_inst.mem.rMemory[6][4] ),
    .A1(_05488_),
    .S(_05601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05606_));
 sky130_fd_sc_hd__clkbuf_1 _12162_ (.A(_05606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00484_));
 sky130_fd_sc_hd__buf_2 _12163_ (.A(_05599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05607_));
 sky130_fd_sc_hd__mux2_1 _12164_ (.A0(\fifo_inst.mem.rMemory[6][5] ),
    .A1(_05490_),
    .S(_05607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05608_));
 sky130_fd_sc_hd__clkbuf_1 _12165_ (.A(_05608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _12166_ (.A0(\fifo_inst.mem.rMemory[6][6] ),
    .A1(_05493_),
    .S(_05607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05609_));
 sky130_fd_sc_hd__clkbuf_1 _12167_ (.A(_05609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _12168_ (.A0(\fifo_inst.mem.rMemory[6][7] ),
    .A1(_05495_),
    .S(_05607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05610_));
 sky130_fd_sc_hd__clkbuf_1 _12169_ (.A(_05610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _12170_ (.A0(\fifo_inst.mem.rMemory[6][8] ),
    .A1(_05497_),
    .S(_05607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05611_));
 sky130_fd_sc_hd__clkbuf_1 _12171_ (.A(_05611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_1 _12172_ (.A0(\fifo_inst.mem.rMemory[6][9] ),
    .A1(_05499_),
    .S(_05607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05612_));
 sky130_fd_sc_hd__clkbuf_1 _12173_ (.A(_05612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00489_));
 sky130_fd_sc_hd__buf_2 _12174_ (.A(_05599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05613_));
 sky130_fd_sc_hd__mux2_1 _12175_ (.A0(\fifo_inst.mem.rMemory[6][10] ),
    .A1(_05501_),
    .S(_05613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05614_));
 sky130_fd_sc_hd__clkbuf_1 _12176_ (.A(_05614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _12177_ (.A0(\fifo_inst.mem.rMemory[6][11] ),
    .A1(_05504_),
    .S(_05613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05615_));
 sky130_fd_sc_hd__clkbuf_1 _12178_ (.A(_05615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _12179_ (.A0(\fifo_inst.mem.rMemory[6][12] ),
    .A1(_05506_),
    .S(_05613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05616_));
 sky130_fd_sc_hd__clkbuf_1 _12180_ (.A(_05616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _12181_ (.A0(\fifo_inst.mem.rMemory[6][13] ),
    .A1(_05508_),
    .S(_05613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05617_));
 sky130_fd_sc_hd__clkbuf_1 _12182_ (.A(_05617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _12183_ (.A0(\fifo_inst.mem.rMemory[6][14] ),
    .A1(_05510_),
    .S(_05613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05618_));
 sky130_fd_sc_hd__clkbuf_1 _12184_ (.A(_05618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00494_));
 sky130_fd_sc_hd__buf_2 _12185_ (.A(_05599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05619_));
 sky130_fd_sc_hd__mux2_1 _12186_ (.A0(\fifo_inst.mem.rMemory[6][15] ),
    .A1(_05512_),
    .S(_05619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05620_));
 sky130_fd_sc_hd__clkbuf_1 _12187_ (.A(_05620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _12188_ (.A0(\fifo_inst.mem.rMemory[6][16] ),
    .A1(_05515_),
    .S(_05619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05621_));
 sky130_fd_sc_hd__clkbuf_1 _12189_ (.A(_05621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_1 _12190_ (.A0(\fifo_inst.mem.rMemory[6][17] ),
    .A1(_05517_),
    .S(_05619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05622_));
 sky130_fd_sc_hd__clkbuf_1 _12191_ (.A(_05622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _12192_ (.A0(\fifo_inst.mem.rMemory[6][18] ),
    .A1(_05519_),
    .S(_05619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05623_));
 sky130_fd_sc_hd__clkbuf_1 _12193_ (.A(_05623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00498_));
 sky130_fd_sc_hd__mux2_1 _12194_ (.A0(\fifo_inst.mem.rMemory[6][19] ),
    .A1(_05521_),
    .S(_05619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05624_));
 sky130_fd_sc_hd__clkbuf_1 _12195_ (.A(_05624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _12196_ (.A0(\fifo_inst.mem.rMemory[6][20] ),
    .A1(_05523_),
    .S(_05600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05625_));
 sky130_fd_sc_hd__clkbuf_1 _12197_ (.A(_05625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _12198_ (.A0(\fifo_inst.mem.rMemory[6][21] ),
    .A1(_05525_),
    .S(_05600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05626_));
 sky130_fd_sc_hd__clkbuf_1 _12199_ (.A(_05626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _12200_ (.A0(\fifo_inst.mem.rMemory[6][22] ),
    .A1(_05527_),
    .S(_05600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05627_));
 sky130_fd_sc_hd__clkbuf_1 _12201_ (.A(_05627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _12202_ (.A0(\fifo_inst.mem.rMemory[6][23] ),
    .A1(_05529_),
    .S(_05600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05628_));
 sky130_fd_sc_hd__clkbuf_1 _12203_ (.A(_05628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00503_));
 sky130_fd_sc_hd__nor2_1 _12204_ (.A(\sa_inst.cols_l2a:2.l2a_i._27_ ),
    .B(\sa_inst.cols_l2a:2.l2a_i._23_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05629_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12205_ (.A(_05629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05630_));
 sky130_fd_sc_hd__o21ai_1 _12206_ (.A1(\sa_inst.cols_l2a:2.l2a_i._09_[0] ),
    .A2(\sa_inst.cols_l2a:2.l2a_i._15_ ),
    .B1(_05630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05631_));
 sky130_fd_sc_hd__a21oi_1 _12207_ (.A1(\sa_inst.cols_l2a:2.l2a_i._09_[0] ),
    .A2(\sa_inst.cols_l2a:2.l2a_i._15_ ),
    .B1(_05631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00504_));
 sky130_fd_sc_hd__and3_1 _12208_ (.A(\sa_inst.cols_l2a:2.l2a_i._09_[0] ),
    .B(\sa_inst.cols_l2a:2.l2a_i._15_ ),
    .C(\sa_inst.cols_l2a:2.l2a_i._09_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05632_));
 sky130_fd_sc_hd__a21o_1 _12209_ (.A1(\sa_inst.cols_l2a:2.l2a_i._09_[0] ),
    .A2(\sa_inst.cols_l2a:2.l2a_i._15_ ),
    .B1(\sa_inst.cols_l2a:2.l2a_i._09_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05633_));
 sky130_fd_sc_hd__and3b_1 _12210_ (.A_N(_05632_),
    .B(_05629_),
    .C(_05633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05634_));
 sky130_fd_sc_hd__clkbuf_1 _12211_ (.A(_05634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00505_));
 sky130_fd_sc_hd__and2_1 _12212_ (.A(\sa_inst.cols_l2a:2.l2a_i._09_[2] ),
    .B(_05632_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05635_));
 sky130_fd_sc_hd__o21ai_1 _12213_ (.A1(\sa_inst.cols_l2a:2.l2a_i._09_[2] ),
    .A2(_05632_),
    .B1(_05630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05636_));
 sky130_fd_sc_hd__nor2_1 _12214_ (.A(_05635_),
    .B(_05636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00506_));
 sky130_fd_sc_hd__and3_1 _12215_ (.A(\sa_inst.cols_l2a:2.l2a_i._09_[2] ),
    .B(\sa_inst.cols_l2a:2.l2a_i._09_[3] ),
    .C(_05632_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05637_));
 sky130_fd_sc_hd__o21ai_1 _12216_ (.A1(\sa_inst.cols_l2a:2.l2a_i._09_[3] ),
    .A2(_05635_),
    .B1(_05630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05638_));
 sky130_fd_sc_hd__nor2_1 _12217_ (.A(_05637_),
    .B(_05638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00507_));
 sky130_fd_sc_hd__o21ai_1 _12218_ (.A1(\sa_inst.cols_l2a:2.l2a_i._09_[4] ),
    .A2(_05637_),
    .B1(_05630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05639_));
 sky130_fd_sc_hd__a21oi_1 _12219_ (.A1(\sa_inst.cols_l2a:2.l2a_i._09_[4] ),
    .A2(_05637_),
    .B1(_05639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00508_));
 sky130_fd_sc_hd__and3_1 _12220_ (.A(\sa_inst.cols_l2a:2.l2a_i._09_[4] ),
    .B(\sa_inst.cols_l2a:2.l2a_i._09_[5] ),
    .C(_05637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05640_));
 sky130_fd_sc_hd__a21o_1 _12221_ (.A1(\sa_inst.cols_l2a:2.l2a_i._09_[4] ),
    .A2(_05637_),
    .B1(\sa_inst.cols_l2a:2.l2a_i._09_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05641_));
 sky130_fd_sc_hd__and3b_1 _12222_ (.A_N(_05640_),
    .B(_05629_),
    .C(_05641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05642_));
 sky130_fd_sc_hd__clkbuf_1 _12223_ (.A(_05642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00509_));
 sky130_fd_sc_hd__a21boi_1 _12224_ (.A1(\sa_inst.cols_l2a:2.l2a_i._09_[6] ),
    .A2(_05640_),
    .B1_N(_05630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05643_));
 sky130_fd_sc_hd__o21a_1 _12225_ (.A1(\sa_inst.cols_l2a:2.l2a_i._09_[6] ),
    .A2(_05640_),
    .B1(_05643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00510_));
 sky130_fd_sc_hd__or2b_4 _12226_ (.A(_05184_),
    .B_N(_05344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05644_));
 sky130_fd_sc_hd__buf_2 _12227_ (.A(_05644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05645_));
 sky130_fd_sc_hd__buf_2 _12228_ (.A(_05645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05646_));
 sky130_fd_sc_hd__mux2_1 _12229_ (.A0(_05064_),
    .A1(\fifo_inst.mem.rMemory[15][0] ),
    .S(_05646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05647_));
 sky130_fd_sc_hd__clkbuf_1 _12230_ (.A(_05647_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _12231_ (.A0(_05076_),
    .A1(\fifo_inst.mem.rMemory[15][1] ),
    .S(_05646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05648_));
 sky130_fd_sc_hd__clkbuf_1 _12232_ (.A(_05648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _12233_ (.A0(_05078_),
    .A1(\fifo_inst.mem.rMemory[15][2] ),
    .S(_05646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05649_));
 sky130_fd_sc_hd__clkbuf_1 _12234_ (.A(_05649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _12235_ (.A0(_05080_),
    .A1(\fifo_inst.mem.rMemory[15][3] ),
    .S(_05646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05650_));
 sky130_fd_sc_hd__clkbuf_1 _12236_ (.A(_05650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _12237_ (.A0(_05082_),
    .A1(\fifo_inst.mem.rMemory[15][4] ),
    .S(_05646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05651_));
 sky130_fd_sc_hd__clkbuf_1 _12238_ (.A(_05651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00515_));
 sky130_fd_sc_hd__buf_2 _12239_ (.A(_05644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05652_));
 sky130_fd_sc_hd__mux2_1 _12240_ (.A0(_05084_),
    .A1(\fifo_inst.mem.rMemory[15][5] ),
    .S(_05652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05653_));
 sky130_fd_sc_hd__clkbuf_1 _12241_ (.A(_05653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _12242_ (.A0(_05087_),
    .A1(\fifo_inst.mem.rMemory[15][6] ),
    .S(_05652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05654_));
 sky130_fd_sc_hd__clkbuf_1 _12243_ (.A(_05654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _12244_ (.A0(_05089_),
    .A1(\fifo_inst.mem.rMemory[15][7] ),
    .S(_05652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05655_));
 sky130_fd_sc_hd__clkbuf_1 _12245_ (.A(_05655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_1 _12246_ (.A0(_05091_),
    .A1(\fifo_inst.mem.rMemory[15][8] ),
    .S(_05652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05656_));
 sky130_fd_sc_hd__clkbuf_1 _12247_ (.A(_05656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _12248_ (.A0(_05093_),
    .A1(\fifo_inst.mem.rMemory[15][9] ),
    .S(_05652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05657_));
 sky130_fd_sc_hd__clkbuf_1 _12249_ (.A(_05657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00520_));
 sky130_fd_sc_hd__buf_2 _12250_ (.A(_05644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05658_));
 sky130_fd_sc_hd__mux2_1 _12251_ (.A0(_05095_),
    .A1(\fifo_inst.mem.rMemory[15][10] ),
    .S(_05658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05659_));
 sky130_fd_sc_hd__clkbuf_1 _12252_ (.A(_05659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _12253_ (.A0(_05098_),
    .A1(\fifo_inst.mem.rMemory[15][11] ),
    .S(_05658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05660_));
 sky130_fd_sc_hd__clkbuf_1 _12254_ (.A(_05660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_1 _12255_ (.A0(_05100_),
    .A1(\fifo_inst.mem.rMemory[15][12] ),
    .S(_05658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05661_));
 sky130_fd_sc_hd__clkbuf_1 _12256_ (.A(_05661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _12257_ (.A0(_05102_),
    .A1(\fifo_inst.mem.rMemory[15][13] ),
    .S(_05658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05662_));
 sky130_fd_sc_hd__clkbuf_1 _12258_ (.A(_05662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _12259_ (.A0(_05104_),
    .A1(\fifo_inst.mem.rMemory[15][14] ),
    .S(_05658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05663_));
 sky130_fd_sc_hd__clkbuf_1 _12260_ (.A(_05663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00525_));
 sky130_fd_sc_hd__buf_2 _12261_ (.A(_05644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05664_));
 sky130_fd_sc_hd__mux2_1 _12262_ (.A0(_05106_),
    .A1(\fifo_inst.mem.rMemory[15][15] ),
    .S(_05664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05665_));
 sky130_fd_sc_hd__clkbuf_1 _12263_ (.A(_05665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _12264_ (.A0(_05113_),
    .A1(\fifo_inst.mem.rMemory[15][16] ),
    .S(_05664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05666_));
 sky130_fd_sc_hd__clkbuf_1 _12265_ (.A(_05666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _12266_ (.A0(_05118_),
    .A1(\fifo_inst.mem.rMemory[15][17] ),
    .S(_05664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05667_));
 sky130_fd_sc_hd__clkbuf_1 _12267_ (.A(_05667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_1 _12268_ (.A0(_05122_),
    .A1(\fifo_inst.mem.rMemory[15][18] ),
    .S(_05664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05668_));
 sky130_fd_sc_hd__clkbuf_1 _12269_ (.A(_05668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _12270_ (.A0(_05127_),
    .A1(\fifo_inst.mem.rMemory[15][19] ),
    .S(_05664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05669_));
 sky130_fd_sc_hd__clkbuf_1 _12271_ (.A(_05669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _12272_ (.A0(_05131_),
    .A1(\fifo_inst.mem.rMemory[15][20] ),
    .S(_05645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05670_));
 sky130_fd_sc_hd__clkbuf_1 _12273_ (.A(_05670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _12274_ (.A0(_05136_),
    .A1(\fifo_inst.mem.rMemory[15][21] ),
    .S(_05645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05671_));
 sky130_fd_sc_hd__clkbuf_1 _12275_ (.A(_05671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _12276_ (.A0(_05140_),
    .A1(\fifo_inst.mem.rMemory[15][22] ),
    .S(_05645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05672_));
 sky130_fd_sc_hd__clkbuf_1 _12277_ (.A(_05672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _12278_ (.A0(_05144_),
    .A1(\fifo_inst.mem.rMemory[15][23] ),
    .S(_05645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05673_));
 sky130_fd_sc_hd__clkbuf_1 _12279_ (.A(_05673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00534_));
 sky130_fd_sc_hd__nor2_4 _12280_ (.A(_05280_),
    .B(_05598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05674_));
 sky130_fd_sc_hd__buf_2 _12281_ (.A(_05674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05675_));
 sky130_fd_sc_hd__buf_2 _12282_ (.A(_05675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05676_));
 sky130_fd_sc_hd__mux2_1 _12283_ (.A0(\fifo_inst.mem.rMemory[5][0] ),
    .A1(_05477_),
    .S(_05676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05677_));
 sky130_fd_sc_hd__clkbuf_1 _12284_ (.A(_05677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _12285_ (.A0(\fifo_inst.mem.rMemory[5][1] ),
    .A1(_05482_),
    .S(_05676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05678_));
 sky130_fd_sc_hd__clkbuf_1 _12286_ (.A(_05678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _12287_ (.A0(\fifo_inst.mem.rMemory[5][2] ),
    .A1(_05484_),
    .S(_05676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05679_));
 sky130_fd_sc_hd__clkbuf_1 _12288_ (.A(_05679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _12289_ (.A0(\fifo_inst.mem.rMemory[5][3] ),
    .A1(_05486_),
    .S(_05676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05680_));
 sky130_fd_sc_hd__clkbuf_1 _12290_ (.A(_05680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_1 _12291_ (.A0(\fifo_inst.mem.rMemory[5][4] ),
    .A1(_05488_),
    .S(_05676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05681_));
 sky130_fd_sc_hd__clkbuf_1 _12292_ (.A(_05681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00539_));
 sky130_fd_sc_hd__buf_2 _12293_ (.A(_05674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05682_));
 sky130_fd_sc_hd__mux2_1 _12294_ (.A0(\fifo_inst.mem.rMemory[5][5] ),
    .A1(_05490_),
    .S(_05682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05683_));
 sky130_fd_sc_hd__clkbuf_1 _12295_ (.A(_05683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_1 _12296_ (.A0(\fifo_inst.mem.rMemory[5][6] ),
    .A1(_05493_),
    .S(_05682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05684_));
 sky130_fd_sc_hd__clkbuf_1 _12297_ (.A(_05684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00541_));
 sky130_fd_sc_hd__mux2_1 _12298_ (.A0(\fifo_inst.mem.rMemory[5][7] ),
    .A1(_05495_),
    .S(_05682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05685_));
 sky130_fd_sc_hd__clkbuf_1 _12299_ (.A(_05685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_1 _12300_ (.A0(\fifo_inst.mem.rMemory[5][8] ),
    .A1(_05497_),
    .S(_05682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05686_));
 sky130_fd_sc_hd__clkbuf_1 _12301_ (.A(_05686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00543_));
 sky130_fd_sc_hd__mux2_1 _12302_ (.A0(\fifo_inst.mem.rMemory[5][9] ),
    .A1(_05499_),
    .S(_05682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05687_));
 sky130_fd_sc_hd__clkbuf_1 _12303_ (.A(_05687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00544_));
 sky130_fd_sc_hd__buf_2 _12304_ (.A(_05674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05688_));
 sky130_fd_sc_hd__mux2_1 _12305_ (.A0(\fifo_inst.mem.rMemory[5][10] ),
    .A1(_05501_),
    .S(_05688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05689_));
 sky130_fd_sc_hd__clkbuf_1 _12306_ (.A(_05689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00545_));
 sky130_fd_sc_hd__mux2_1 _12307_ (.A0(\fifo_inst.mem.rMemory[5][11] ),
    .A1(_05504_),
    .S(_05688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05690_));
 sky130_fd_sc_hd__clkbuf_1 _12308_ (.A(_05690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_1 _12309_ (.A0(\fifo_inst.mem.rMemory[5][12] ),
    .A1(_05506_),
    .S(_05688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05691_));
 sky130_fd_sc_hd__clkbuf_1 _12310_ (.A(_05691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _12311_ (.A0(\fifo_inst.mem.rMemory[5][13] ),
    .A1(_05508_),
    .S(_05688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05692_));
 sky130_fd_sc_hd__clkbuf_1 _12312_ (.A(_05692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_1 _12313_ (.A0(\fifo_inst.mem.rMemory[5][14] ),
    .A1(_05510_),
    .S(_05688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05693_));
 sky130_fd_sc_hd__clkbuf_1 _12314_ (.A(_05693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00549_));
 sky130_fd_sc_hd__buf_2 _12315_ (.A(_05674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05694_));
 sky130_fd_sc_hd__mux2_1 _12316_ (.A0(\fifo_inst.mem.rMemory[5][15] ),
    .A1(_05512_),
    .S(_05694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05695_));
 sky130_fd_sc_hd__clkbuf_1 _12317_ (.A(_05695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _12318_ (.A0(\fifo_inst.mem.rMemory[5][16] ),
    .A1(_05515_),
    .S(_05694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05696_));
 sky130_fd_sc_hd__clkbuf_1 _12319_ (.A(_05696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _12320_ (.A0(\fifo_inst.mem.rMemory[5][17] ),
    .A1(_05517_),
    .S(_05694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05697_));
 sky130_fd_sc_hd__clkbuf_1 _12321_ (.A(_05697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _12322_ (.A0(\fifo_inst.mem.rMemory[5][18] ),
    .A1(_05519_),
    .S(_05694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05698_));
 sky130_fd_sc_hd__clkbuf_1 _12323_ (.A(_05698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_1 _12324_ (.A0(\fifo_inst.mem.rMemory[5][19] ),
    .A1(_05521_),
    .S(_05694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05699_));
 sky130_fd_sc_hd__clkbuf_1 _12325_ (.A(_05699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _12326_ (.A0(\fifo_inst.mem.rMemory[5][20] ),
    .A1(_05523_),
    .S(_05675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05700_));
 sky130_fd_sc_hd__clkbuf_1 _12327_ (.A(_05700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _12328_ (.A0(\fifo_inst.mem.rMemory[5][21] ),
    .A1(_05525_),
    .S(_05675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05701_));
 sky130_fd_sc_hd__clkbuf_1 _12329_ (.A(_05701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _12330_ (.A0(\fifo_inst.mem.rMemory[5][22] ),
    .A1(_05527_),
    .S(_05675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05702_));
 sky130_fd_sc_hd__clkbuf_1 _12331_ (.A(_05702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _12332_ (.A0(\fifo_inst.mem.rMemory[5][23] ),
    .A1(_05529_),
    .S(_05675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05703_));
 sky130_fd_sc_hd__clkbuf_1 _12333_ (.A(_05703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00558_));
 sky130_fd_sc_hd__and3_1 _12334_ (.A(\sa_inst._00_[0] ),
    .B(_01037_),
    .C(_00810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05704_));
 sky130_fd_sc_hd__clkbuf_1 _12335_ (.A(_05704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00559_));
 sky130_fd_sc_hd__and3_1 _12336_ (.A(\sa_inst._00_[1] ),
    .B(_01037_),
    .C(_00810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05705_));
 sky130_fd_sc_hd__clkbuf_1 _12337_ (.A(_05705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00560_));
 sky130_fd_sc_hd__and2_1 _12338_ (.A(\sa_inst._00_[2] ),
    .B(_01037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05706_));
 sky130_fd_sc_hd__clkbuf_1 _12339_ (.A(_05706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00561_));
 sky130_fd_sc_hd__and2_1 _12340_ (.A(\sa_inst._00_[3] ),
    .B(_01037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05707_));
 sky130_fd_sc_hd__clkbuf_1 _12341_ (.A(_05707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00562_));
 sky130_fd_sc_hd__nor2_4 _12342_ (.A(_05311_),
    .B(_05598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05708_));
 sky130_fd_sc_hd__buf_2 _12343_ (.A(_05708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05709_));
 sky130_fd_sc_hd__buf_2 _12344_ (.A(_05709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05710_));
 sky130_fd_sc_hd__mux2_1 _12345_ (.A0(\fifo_inst.mem.rMemory[4][0] ),
    .A1(_05477_),
    .S(_05710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05711_));
 sky130_fd_sc_hd__clkbuf_1 _12346_ (.A(_05711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _12347_ (.A0(\fifo_inst.mem.rMemory[4][1] ),
    .A1(_05482_),
    .S(_05710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05712_));
 sky130_fd_sc_hd__clkbuf_1 _12348_ (.A(_05712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _12349_ (.A0(\fifo_inst.mem.rMemory[4][2] ),
    .A1(_05484_),
    .S(_05710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05713_));
 sky130_fd_sc_hd__clkbuf_1 _12350_ (.A(_05713_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _12351_ (.A0(\fifo_inst.mem.rMemory[4][3] ),
    .A1(_05486_),
    .S(_05710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05714_));
 sky130_fd_sc_hd__clkbuf_1 _12352_ (.A(_05714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_1 _12353_ (.A0(\fifo_inst.mem.rMemory[4][4] ),
    .A1(_05488_),
    .S(_05710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05715_));
 sky130_fd_sc_hd__clkbuf_1 _12354_ (.A(_05715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00567_));
 sky130_fd_sc_hd__buf_2 _12355_ (.A(_05708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05716_));
 sky130_fd_sc_hd__mux2_1 _12356_ (.A0(\fifo_inst.mem.rMemory[4][5] ),
    .A1(_05490_),
    .S(_05716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05717_));
 sky130_fd_sc_hd__clkbuf_1 _12357_ (.A(_05717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _12358_ (.A0(\fifo_inst.mem.rMemory[4][6] ),
    .A1(_05493_),
    .S(_05716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05718_));
 sky130_fd_sc_hd__clkbuf_1 _12359_ (.A(_05718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _12360_ (.A0(\fifo_inst.mem.rMemory[4][7] ),
    .A1(_05495_),
    .S(_05716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05719_));
 sky130_fd_sc_hd__clkbuf_1 _12361_ (.A(_05719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _12362_ (.A0(\fifo_inst.mem.rMemory[4][8] ),
    .A1(_05497_),
    .S(_05716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05720_));
 sky130_fd_sc_hd__clkbuf_1 _12363_ (.A(_05720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _12364_ (.A0(\fifo_inst.mem.rMemory[4][9] ),
    .A1(_05499_),
    .S(_05716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05721_));
 sky130_fd_sc_hd__clkbuf_1 _12365_ (.A(_05721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00572_));
 sky130_fd_sc_hd__buf_2 _12366_ (.A(_05708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05722_));
 sky130_fd_sc_hd__mux2_1 _12367_ (.A0(\fifo_inst.mem.rMemory[4][10] ),
    .A1(_05501_),
    .S(_05722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05723_));
 sky130_fd_sc_hd__clkbuf_1 _12368_ (.A(_05723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_1 _12369_ (.A0(\fifo_inst.mem.rMemory[4][11] ),
    .A1(_05504_),
    .S(_05722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05724_));
 sky130_fd_sc_hd__clkbuf_1 _12370_ (.A(_05724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_1 _12371_ (.A0(\fifo_inst.mem.rMemory[4][12] ),
    .A1(_05506_),
    .S(_05722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05725_));
 sky130_fd_sc_hd__clkbuf_1 _12372_ (.A(_05725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _12373_ (.A0(\fifo_inst.mem.rMemory[4][13] ),
    .A1(_05508_),
    .S(_05722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05726_));
 sky130_fd_sc_hd__clkbuf_1 _12374_ (.A(_05726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _12375_ (.A0(\fifo_inst.mem.rMemory[4][14] ),
    .A1(_05510_),
    .S(_05722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05727_));
 sky130_fd_sc_hd__clkbuf_1 _12376_ (.A(_05727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00577_));
 sky130_fd_sc_hd__buf_2 _12377_ (.A(_05708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05728_));
 sky130_fd_sc_hd__mux2_1 _12378_ (.A0(\fifo_inst.mem.rMemory[4][15] ),
    .A1(_05512_),
    .S(_05728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05729_));
 sky130_fd_sc_hd__clkbuf_1 _12379_ (.A(_05729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _12380_ (.A0(\fifo_inst.mem.rMemory[4][16] ),
    .A1(_05515_),
    .S(_05728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05730_));
 sky130_fd_sc_hd__clkbuf_1 _12381_ (.A(_05730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _12382_ (.A0(\fifo_inst.mem.rMemory[4][17] ),
    .A1(_05517_),
    .S(_05728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05731_));
 sky130_fd_sc_hd__clkbuf_1 _12383_ (.A(_05731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _12384_ (.A0(\fifo_inst.mem.rMemory[4][18] ),
    .A1(_05519_),
    .S(_05728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05732_));
 sky130_fd_sc_hd__clkbuf_1 _12385_ (.A(_05732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _12386_ (.A0(\fifo_inst.mem.rMemory[4][19] ),
    .A1(_05521_),
    .S(_05728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05733_));
 sky130_fd_sc_hd__clkbuf_1 _12387_ (.A(_05733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _12388_ (.A0(\fifo_inst.mem.rMemory[4][20] ),
    .A1(_05523_),
    .S(_05709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05734_));
 sky130_fd_sc_hd__clkbuf_1 _12389_ (.A(_05734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _12390_ (.A0(\fifo_inst.mem.rMemory[4][21] ),
    .A1(_05525_),
    .S(_05709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05735_));
 sky130_fd_sc_hd__clkbuf_1 _12391_ (.A(_05735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _12392_ (.A0(\fifo_inst.mem.rMemory[4][22] ),
    .A1(_05527_),
    .S(_05709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05736_));
 sky130_fd_sc_hd__clkbuf_1 _12393_ (.A(_05736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _12394_ (.A0(\fifo_inst.mem.rMemory[4][23] ),
    .A1(_05529_),
    .S(_05709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05737_));
 sky130_fd_sc_hd__clkbuf_1 _12395_ (.A(_05737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00586_));
 sky130_fd_sc_hd__and3_1 _12396_ (.A(net1),
    .B(_04315_),
    .C(_00820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05738_));
 sky130_fd_sc_hd__clkbuf_1 _12397_ (.A(_05738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00587_));
 sky130_fd_sc_hd__and3_1 _12398_ (.A(net12),
    .B(_04315_),
    .C(_00820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05739_));
 sky130_fd_sc_hd__clkbuf_1 _12399_ (.A(_05739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00588_));
 sky130_fd_sc_hd__and3_1 _12400_ (.A(net17),
    .B(_04315_),
    .C(_00820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05740_));
 sky130_fd_sc_hd__clkbuf_1 _12401_ (.A(_05740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00589_));
 sky130_fd_sc_hd__and3b_1 _12402_ (.A_N(_00819_),
    .B(_04315_),
    .C(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05741_));
 sky130_fd_sc_hd__clkbuf_1 _12403_ (.A(_05741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00590_));
 sky130_fd_sc_hd__and2b_1 _12404_ (.A_N(_04125_),
    .B(_04122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05742_));
 sky130_fd_sc_hd__clkbuf_1 _12405_ (.A(_05742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00591_));
 sky130_fd_sc_hd__buf_2 _12406_ (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05743_));
 sky130_fd_sc_hd__clkbuf_1 _12407_ (.A(_05743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05744_));
 sky130_fd_sc_hd__buf_2 _12408_ (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05745_));
 sky130_fd_sc_hd__clkbuf_1 _12409_ (.A(_05745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05746_));
 sky130_fd_sc_hd__and3_1 _12410_ (.A(_05744_),
    .B(_05746_),
    .C(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05747_));
 sky130_fd_sc_hd__clkbuf_1 _12411_ (.A(_05747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00592_));
 sky130_fd_sc_hd__and3_1 _12412_ (.A(_05744_),
    .B(_05746_),
    .C(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05748_));
 sky130_fd_sc_hd__clkbuf_1 _12413_ (.A(_05748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00593_));
 sky130_fd_sc_hd__and3_1 _12414_ (.A(_05744_),
    .B(_05746_),
    .C(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05749_));
 sky130_fd_sc_hd__clkbuf_1 _12415_ (.A(_05749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00594_));
 sky130_fd_sc_hd__and3_1 _12416_ (.A(_05744_),
    .B(_05746_),
    .C(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05750_));
 sky130_fd_sc_hd__clkbuf_1 _12417_ (.A(_05750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00595_));
 sky130_fd_sc_hd__and3_1 _12418_ (.A(_05744_),
    .B(_05746_),
    .C(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05751_));
 sky130_fd_sc_hd__clkbuf_1 _12419_ (.A(_05751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00596_));
 sky130_fd_sc_hd__clkbuf_1 _12420_ (.A(_05743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05752_));
 sky130_fd_sc_hd__clkbuf_1 _12421_ (.A(_05745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05753_));
 sky130_fd_sc_hd__and3_1 _12422_ (.A(_05752_),
    .B(_05753_),
    .C(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05754_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12423_ (.A(_05754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00597_));
 sky130_fd_sc_hd__and3_1 _12424_ (.A(_05752_),
    .B(_05753_),
    .C(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05755_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12425_ (.A(_05755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00598_));
 sky130_fd_sc_hd__and3_1 _12426_ (.A(_05752_),
    .B(_05753_),
    .C(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05756_));
 sky130_fd_sc_hd__clkbuf_1 _12427_ (.A(_05756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00599_));
 sky130_fd_sc_hd__nor2_8 _12428_ (.A(_05071_),
    .B(_05280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05757_));
 sky130_fd_sc_hd__buf_2 _12429_ (.A(_05757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05758_));
 sky130_fd_sc_hd__buf_2 _12430_ (.A(_05758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05759_));
 sky130_fd_sc_hd__mux2_1 _12431_ (.A0(\fifo_inst.mem.rMemory[1][0] ),
    .A1(\fifo_inst.WR_DATA[0] ),
    .S(_05759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05760_));
 sky130_fd_sc_hd__clkbuf_1 _12432_ (.A(_05760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _12433_ (.A0(\fifo_inst.mem.rMemory[1][1] ),
    .A1(\fifo_inst.WR_DATA[1] ),
    .S(_05759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05761_));
 sky130_fd_sc_hd__clkbuf_1 _12434_ (.A(_05761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _12435_ (.A0(\fifo_inst.mem.rMemory[1][2] ),
    .A1(\fifo_inst.WR_DATA[2] ),
    .S(_05759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05762_));
 sky130_fd_sc_hd__clkbuf_1 _12436_ (.A(_05762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _12437_ (.A0(\fifo_inst.mem.rMemory[1][3] ),
    .A1(\fifo_inst.WR_DATA[3] ),
    .S(_05759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05763_));
 sky130_fd_sc_hd__clkbuf_1 _12438_ (.A(_05763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _12439_ (.A0(\fifo_inst.mem.rMemory[1][4] ),
    .A1(\fifo_inst.WR_DATA[4] ),
    .S(_05759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05764_));
 sky130_fd_sc_hd__clkbuf_1 _12440_ (.A(_05764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00604_));
 sky130_fd_sc_hd__buf_2 _12441_ (.A(_05757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05765_));
 sky130_fd_sc_hd__mux2_1 _12442_ (.A0(\fifo_inst.mem.rMemory[1][5] ),
    .A1(\fifo_inst.WR_DATA[5] ),
    .S(_05765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05766_));
 sky130_fd_sc_hd__clkbuf_1 _12443_ (.A(_05766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _12444_ (.A0(\fifo_inst.mem.rMemory[1][6] ),
    .A1(\fifo_inst.WR_DATA[6] ),
    .S(_05765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05767_));
 sky130_fd_sc_hd__clkbuf_1 _12445_ (.A(_05767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _12446_ (.A0(\fifo_inst.mem.rMemory[1][7] ),
    .A1(\fifo_inst.WR_DATA[7] ),
    .S(_05765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05768_));
 sky130_fd_sc_hd__clkbuf_1 _12447_ (.A(_05768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _12448_ (.A0(\fifo_inst.mem.rMemory[1][8] ),
    .A1(\fifo_inst.WR_DATA[8] ),
    .S(_05765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05769_));
 sky130_fd_sc_hd__clkbuf_1 _12449_ (.A(_05769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_1 _12450_ (.A0(\fifo_inst.mem.rMemory[1][9] ),
    .A1(\fifo_inst.WR_DATA[9] ),
    .S(_05765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05770_));
 sky130_fd_sc_hd__clkbuf_1 _12451_ (.A(_05770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00609_));
 sky130_fd_sc_hd__buf_2 _12452_ (.A(_05757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05771_));
 sky130_fd_sc_hd__mux2_1 _12453_ (.A0(\fifo_inst.mem.rMemory[1][10] ),
    .A1(\fifo_inst.WR_DATA[10] ),
    .S(_05771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05772_));
 sky130_fd_sc_hd__clkbuf_1 _12454_ (.A(_05772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _12455_ (.A0(\fifo_inst.mem.rMemory[1][11] ),
    .A1(\fifo_inst.WR_DATA[11] ),
    .S(_05771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05773_));
 sky130_fd_sc_hd__clkbuf_1 _12456_ (.A(_05773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _12457_ (.A0(\fifo_inst.mem.rMemory[1][12] ),
    .A1(\fifo_inst.WR_DATA[12] ),
    .S(_05771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05774_));
 sky130_fd_sc_hd__clkbuf_1 _12458_ (.A(_05774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _12459_ (.A0(\fifo_inst.mem.rMemory[1][13] ),
    .A1(\fifo_inst.WR_DATA[13] ),
    .S(_05771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05775_));
 sky130_fd_sc_hd__clkbuf_1 _12460_ (.A(_05775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_1 _12461_ (.A0(\fifo_inst.mem.rMemory[1][14] ),
    .A1(\fifo_inst.WR_DATA[14] ),
    .S(_05771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05776_));
 sky130_fd_sc_hd__clkbuf_1 _12462_ (.A(_05776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00614_));
 sky130_fd_sc_hd__buf_2 _12463_ (.A(_05757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05777_));
 sky130_fd_sc_hd__mux2_1 _12464_ (.A0(\fifo_inst.mem.rMemory[1][15] ),
    .A1(\fifo_inst.WR_DATA[15] ),
    .S(_05777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05778_));
 sky130_fd_sc_hd__clkbuf_1 _12465_ (.A(_05778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _12466_ (.A0(\fifo_inst.mem.rMemory[1][16] ),
    .A1(_05112_),
    .S(_05777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05779_));
 sky130_fd_sc_hd__clkbuf_1 _12467_ (.A(_05779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_1 _12468_ (.A0(\fifo_inst.mem.rMemory[1][17] ),
    .A1(_05117_),
    .S(_05777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05780_));
 sky130_fd_sc_hd__clkbuf_1 _12469_ (.A(_05780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _12470_ (.A0(\fifo_inst.mem.rMemory[1][18] ),
    .A1(_05121_),
    .S(_05777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05781_));
 sky130_fd_sc_hd__clkbuf_1 _12471_ (.A(_05781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _12472_ (.A0(\fifo_inst.mem.rMemory[1][19] ),
    .A1(_05126_),
    .S(_05777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05782_));
 sky130_fd_sc_hd__clkbuf_1 _12473_ (.A(_05782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _12474_ (.A0(\fifo_inst.mem.rMemory[1][20] ),
    .A1(_05130_),
    .S(_05758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05783_));
 sky130_fd_sc_hd__clkbuf_1 _12475_ (.A(_05783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _12476_ (.A0(\fifo_inst.mem.rMemory[1][21] ),
    .A1(_05135_),
    .S(_05758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05784_));
 sky130_fd_sc_hd__clkbuf_1 _12477_ (.A(_05784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _12478_ (.A0(\fifo_inst.mem.rMemory[1][22] ),
    .A1(_05139_),
    .S(_05758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05785_));
 sky130_fd_sc_hd__clkbuf_1 _12479_ (.A(_05785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _12480_ (.A0(\fifo_inst.mem.rMemory[1][23] ),
    .A1(_05143_),
    .S(_05758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05786_));
 sky130_fd_sc_hd__clkbuf_1 _12481_ (.A(_05786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00623_));
 sky130_fd_sc_hd__and3_1 _12482_ (.A(_05752_),
    .B(_05753_),
    .C(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05787_));
 sky130_fd_sc_hd__clkbuf_1 _12483_ (.A(_05787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00624_));
 sky130_fd_sc_hd__and3_1 _12484_ (.A(_05752_),
    .B(_05753_),
    .C(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05788_));
 sky130_fd_sc_hd__clkbuf_1 _12485_ (.A(_05788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00625_));
 sky130_fd_sc_hd__clkbuf_2 _12486_ (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05789_));
 sky130_fd_sc_hd__clkbuf_2 _12487_ (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05790_));
 sky130_fd_sc_hd__and3_1 _12488_ (.A(_05789_),
    .B(_05790_),
    .C(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05791_));
 sky130_fd_sc_hd__clkbuf_1 _12489_ (.A(_05791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00626_));
 sky130_fd_sc_hd__and3_1 _12490_ (.A(_05789_),
    .B(_05790_),
    .C(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05792_));
 sky130_fd_sc_hd__clkbuf_1 _12491_ (.A(_05792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00627_));
 sky130_fd_sc_hd__and3_1 _12492_ (.A(_05789_),
    .B(_05790_),
    .C(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05793_));
 sky130_fd_sc_hd__clkbuf_1 _12493_ (.A(_05793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00628_));
 sky130_fd_sc_hd__and3_1 _12494_ (.A(_05789_),
    .B(_05790_),
    .C(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05794_));
 sky130_fd_sc_hd__clkbuf_1 _12495_ (.A(_05794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00629_));
 sky130_fd_sc_hd__and3_1 _12496_ (.A(_05789_),
    .B(_05790_),
    .C(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05795_));
 sky130_fd_sc_hd__clkbuf_1 _12497_ (.A(_05795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00630_));
 sky130_fd_sc_hd__and3_1 _12498_ (.A(_05743_),
    .B(_05745_),
    .C(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05796_));
 sky130_fd_sc_hd__clkbuf_1 _12499_ (.A(_05796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00631_));
 sky130_fd_sc_hd__and3_1 _12500_ (.A(_05743_),
    .B(_05745_),
    .C(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05797_));
 sky130_fd_sc_hd__clkbuf_1 _12501_ (.A(_05797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00632_));
 sky130_fd_sc_hd__and3_1 _12502_ (.A(_05743_),
    .B(_05745_),
    .C(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05798_));
 sky130_fd_sc_hd__clkbuf_1 _12503_ (.A(_05798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00633_));
 sky130_fd_sc_hd__inv_2 _12504_ (.A(\sa_inst.cols_l2a:1.l2a_i._27_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05799_));
 sky130_fd_sc_hd__a21o_1 _12505_ (.A1(_05799_),
    .A2(\sa_inst.cols_l2a:1.l2a_i._55_ ),
    .B1(\sa_inst.cols_l2a:1.l2a_i._23_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00634_));
 sky130_fd_sc_hd__inv_2 _12506_ (.A(\sa_inst.cols_l2a:2.l2a_i._27_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05800_));
 sky130_fd_sc_hd__a21o_1 _12507_ (.A1(_05800_),
    .A2(\sa_inst.cols_l2a:2.l2a_i._55_ ),
    .B1(\sa_inst.cols_l2a:2.l2a_i._23_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00635_));
 sky130_fd_sc_hd__and2b_1 _12508_ (.A_N(_04307_),
    .B(_04304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05801_));
 sky130_fd_sc_hd__clkbuf_1 _12509_ (.A(_05801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00636_));
 sky130_fd_sc_hd__or2b_4 _12510_ (.A(_05071_),
    .B_N(_05344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05802_));
 sky130_fd_sc_hd__buf_2 _12511_ (.A(_05802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05803_));
 sky130_fd_sc_hd__buf_2 _12512_ (.A(_05803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05804_));
 sky130_fd_sc_hd__mux2_1 _12513_ (.A0(_05064_),
    .A1(\fifo_inst.mem.rMemory[3][0] ),
    .S(_05804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05805_));
 sky130_fd_sc_hd__clkbuf_1 _12514_ (.A(_05805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _12515_ (.A0(_05076_),
    .A1(\fifo_inst.mem.rMemory[3][1] ),
    .S(_05804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05806_));
 sky130_fd_sc_hd__clkbuf_1 _12516_ (.A(_05806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _12517_ (.A0(_05078_),
    .A1(\fifo_inst.mem.rMemory[3][2] ),
    .S(_05804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05807_));
 sky130_fd_sc_hd__clkbuf_1 _12518_ (.A(_05807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _12519_ (.A0(_05080_),
    .A1(\fifo_inst.mem.rMemory[3][3] ),
    .S(_05804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05808_));
 sky130_fd_sc_hd__clkbuf_1 _12520_ (.A(_05808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _12521_ (.A0(_05082_),
    .A1(\fifo_inst.mem.rMemory[3][4] ),
    .S(_05804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05809_));
 sky130_fd_sc_hd__clkbuf_1 _12522_ (.A(_05809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00641_));
 sky130_fd_sc_hd__buf_2 _12523_ (.A(_05802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05810_));
 sky130_fd_sc_hd__mux2_1 _12524_ (.A0(_05084_),
    .A1(\fifo_inst.mem.rMemory[3][5] ),
    .S(_05810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05811_));
 sky130_fd_sc_hd__clkbuf_1 _12525_ (.A(_05811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _12526_ (.A0(_05087_),
    .A1(\fifo_inst.mem.rMemory[3][6] ),
    .S(_05810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05812_));
 sky130_fd_sc_hd__clkbuf_1 _12527_ (.A(_05812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _12528_ (.A0(_05089_),
    .A1(\fifo_inst.mem.rMemory[3][7] ),
    .S(_05810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05813_));
 sky130_fd_sc_hd__clkbuf_1 _12529_ (.A(_05813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _12530_ (.A0(_05091_),
    .A1(\fifo_inst.mem.rMemory[3][8] ),
    .S(_05810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05814_));
 sky130_fd_sc_hd__clkbuf_1 _12531_ (.A(_05814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _12532_ (.A0(_05093_),
    .A1(\fifo_inst.mem.rMemory[3][9] ),
    .S(_05810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05815_));
 sky130_fd_sc_hd__clkbuf_1 _12533_ (.A(_05815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00646_));
 sky130_fd_sc_hd__buf_2 _12534_ (.A(_05802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05816_));
 sky130_fd_sc_hd__mux2_1 _12535_ (.A0(_05095_),
    .A1(\fifo_inst.mem.rMemory[3][10] ),
    .S(_05816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05817_));
 sky130_fd_sc_hd__clkbuf_1 _12536_ (.A(_05817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _12537_ (.A0(_05098_),
    .A1(\fifo_inst.mem.rMemory[3][11] ),
    .S(_05816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05818_));
 sky130_fd_sc_hd__clkbuf_1 _12538_ (.A(_05818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _12539_ (.A0(_05100_),
    .A1(\fifo_inst.mem.rMemory[3][12] ),
    .S(_05816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05819_));
 sky130_fd_sc_hd__clkbuf_1 _12540_ (.A(_05819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _12541_ (.A0(_05102_),
    .A1(\fifo_inst.mem.rMemory[3][13] ),
    .S(_05816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05820_));
 sky130_fd_sc_hd__clkbuf_1 _12542_ (.A(_05820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _12543_ (.A0(_05104_),
    .A1(\fifo_inst.mem.rMemory[3][14] ),
    .S(_05816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05821_));
 sky130_fd_sc_hd__clkbuf_1 _12544_ (.A(_05821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00651_));
 sky130_fd_sc_hd__buf_2 _12545_ (.A(_05802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05822_));
 sky130_fd_sc_hd__mux2_1 _12546_ (.A0(_05106_),
    .A1(\fifo_inst.mem.rMemory[3][15] ),
    .S(_05822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05823_));
 sky130_fd_sc_hd__clkbuf_1 _12547_ (.A(_05823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _12548_ (.A0(_05113_),
    .A1(\fifo_inst.mem.rMemory[3][16] ),
    .S(_05822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05824_));
 sky130_fd_sc_hd__clkbuf_1 _12549_ (.A(_05824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _12550_ (.A0(_05118_),
    .A1(\fifo_inst.mem.rMemory[3][17] ),
    .S(_05822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05825_));
 sky130_fd_sc_hd__clkbuf_1 _12551_ (.A(_05825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _12552_ (.A0(_05122_),
    .A1(\fifo_inst.mem.rMemory[3][18] ),
    .S(_05822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05826_));
 sky130_fd_sc_hd__clkbuf_1 _12553_ (.A(_05826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _12554_ (.A0(_05127_),
    .A1(\fifo_inst.mem.rMemory[3][19] ),
    .S(_05822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05827_));
 sky130_fd_sc_hd__clkbuf_1 _12555_ (.A(_05827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _12556_ (.A0(_05131_),
    .A1(\fifo_inst.mem.rMemory[3][20] ),
    .S(_05803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05828_));
 sky130_fd_sc_hd__clkbuf_1 _12557_ (.A(_05828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _12558_ (.A0(_05136_),
    .A1(\fifo_inst.mem.rMemory[3][21] ),
    .S(_05803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05829_));
 sky130_fd_sc_hd__clkbuf_1 _12559_ (.A(_05829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _12560_ (.A0(_05140_),
    .A1(\fifo_inst.mem.rMemory[3][22] ),
    .S(_05803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05830_));
 sky130_fd_sc_hd__clkbuf_1 _12561_ (.A(_05830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _12562_ (.A0(_05144_),
    .A1(\fifo_inst.mem.rMemory[3][23] ),
    .S(_05803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05831_));
 sky130_fd_sc_hd__clkbuf_1 _12563_ (.A(_05831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00660_));
 sky130_fd_sc_hd__clkbuf_2 _12564_ (.A(_05343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05832_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12565_ (.A(_05832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05833_));
 sky130_fd_sc_hd__inv_2 _12566_ (.A(_04723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05834_));
 sky130_fd_sc_hd__clkbuf_2 _12567_ (.A(_05834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05835_));
 sky130_fd_sc_hd__inv_2 _12568_ (.A(\fifo_inst.rRdPtrPlus1[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05836_));
 sky130_fd_sc_hd__inv_2 _12569_ (.A(\fifo_inst.rRdPtrPlus1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05837_));
 sky130_fd_sc_hd__inv_2 _12570_ (.A(\fifo_inst.rRdPtrPlus1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05838_));
 sky130_fd_sc_hd__o2bb2a_1 _12571_ (.A1_N(_05837_),
    .A2_N(_05345_),
    .B1(_05342_),
    .B2(_05838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05839_));
 sky130_fd_sc_hd__o221ai_1 _12572_ (.A1(_05836_),
    .A2(\fifo_inst.rWrPtr[4] ),
    .B1(_05345_),
    .B2(_05837_),
    .C1(_05839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05840_));
 sky130_fd_sc_hd__inv_2 _12573_ (.A(\fifo_inst.rRdPtrPlus1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05841_));
 sky130_fd_sc_hd__inv_2 _12574_ (.A(\fifo_inst.rRdPtrPlus1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05842_));
 sky130_fd_sc_hd__a2bb2o_1 _12575_ (.A1_N(_05841_),
    .A2_N(_05278_),
    .B1(\fifo_inst.rWrPtr[4] ),
    .B2(_05836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05843_));
 sky130_fd_sc_hd__a221o_1 _12576_ (.A1(_05838_),
    .A2(_05342_),
    .B1(_05279_),
    .B2(\fifo_inst.rRdPtrPlus1[0] ),
    .C1(_05843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05844_));
 sky130_fd_sc_hd__a221o_1 _12577_ (.A1(_05841_),
    .A2(_05278_),
    .B1(_05065_),
    .B2(_05842_),
    .C1(_05844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05845_));
 sky130_fd_sc_hd__o31a_1 _12578_ (.A1(_05835_),
    .A2(_05840_),
    .A3(_05845_),
    .B1(_04720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05846_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12579_ (.A(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05847_));
 sky130_fd_sc_hd__clkbuf_2 _12580_ (.A(_05847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05848_));
 sky130_fd_sc_hd__o21ai_1 _12581_ (.A1(_05833_),
    .A2(_05846_),
    .B1(_05848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00661_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12582_ (.A(_05067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05849_));
 sky130_fd_sc_hd__or2_1 _12583_ (.A(\fifo_inst.mem.RD1_ADDR[1] ),
    .B(\fifo_inst.rWrPtrPlus1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05850_));
 sky130_fd_sc_hd__nand2_1 _12584_ (.A(_04734_),
    .B(\fifo_inst.rWrPtrPlus1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05851_));
 sky130_fd_sc_hd__or2_1 _12585_ (.A(_04752_),
    .B(\fifo_inst.rWrPtrPlus1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05852_));
 sky130_fd_sc_hd__nand2_1 _12586_ (.A(_04731_),
    .B(\fifo_inst.rWrPtrPlus1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05853_));
 sky130_fd_sc_hd__xor2_1 _12587_ (.A(\fifo_inst.mem.RD1_ADDR[3] ),
    .B(\fifo_inst.rWrPtrPlus1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05854_));
 sky130_fd_sc_hd__a221o_1 _12588_ (.A1(_05850_),
    .A2(_05851_),
    .B1(_05852_),
    .B2(_05853_),
    .C1(_05854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05855_));
 sky130_fd_sc_hd__xnor2_1 _12589_ (.A(\fifo_inst.rRdPtr[4] ),
    .B(\fifo_inst.rWrPtrPlus1[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05856_));
 sky130_fd_sc_hd__xor2_1 _12590_ (.A(_04727_),
    .B(\fifo_inst.rWrPtrPlus1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05857_));
 sky130_fd_sc_hd__or4_1 _12591_ (.A(_05849_),
    .B(_05855_),
    .C(_05856_),
    .D(_05857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05858_));
 sky130_fd_sc_hd__o22a_1 _12592_ (.A1(_04718_),
    .A2(_04719_),
    .B1(_04724_),
    .B2(_05858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05859_));
 sky130_fd_sc_hd__clkbuf_2 _12593_ (.A(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05860_));
 sky130_fd_sc_hd__and2b_1 _12594_ (.A_N(_05859_),
    .B(_05860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05861_));
 sky130_fd_sc_hd__clkbuf_1 _12595_ (.A(_05861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00662_));
 sky130_fd_sc_hd__and2_1 _12596_ (.A(net55),
    .B(_04721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05862_));
 sky130_fd_sc_hd__o21a_1 _12597_ (.A1(_04720_),
    .A2(_05862_),
    .B1(_05848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00663_));
 sky130_fd_sc_hd__and2_1 _12598_ (.A(\fifo_inst.rWrPtrPlus1[0] ),
    .B(_05832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05863_));
 sky130_fd_sc_hd__nor2_1 _12599_ (.A(\fifo_inst.rWrPtrPlus1[0] ),
    .B(_05833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05864_));
 sky130_fd_sc_hd__o21ai_1 _12600_ (.A1(_05863_),
    .A2(_05864_),
    .B1(_05848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00664_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12601_ (.A(\fifo_inst.rWrPtrPlus1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05865_));
 sky130_fd_sc_hd__o21ai_1 _12602_ (.A1(_05865_),
    .A2(_05863_),
    .B1(_05847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05866_));
 sky130_fd_sc_hd__a21oi_1 _12603_ (.A1(_05865_),
    .A2(_05863_),
    .B1(_05866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00665_));
 sky130_fd_sc_hd__and3_1 _12604_ (.A(\fifo_inst.rWrPtrPlus1[2] ),
    .B(_05865_),
    .C(_05863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05867_));
 sky130_fd_sc_hd__a31o_1 _12605_ (.A1(_05865_),
    .A2(\fifo_inst.rWrPtrPlus1[0] ),
    .A3(_05832_),
    .B1(\fifo_inst.rWrPtrPlus1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05868_));
 sky130_fd_sc_hd__and3b_1 _12606_ (.A_N(_05867_),
    .B(_05860_),
    .C(_05868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05869_));
 sky130_fd_sc_hd__clkbuf_1 _12607_ (.A(_05869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00666_));
 sky130_fd_sc_hd__and2_1 _12608_ (.A(\fifo_inst.rWrPtrPlus1[3] ),
    .B(_05867_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05870_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12609_ (.A(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05871_));
 sky130_fd_sc_hd__o21ai_1 _12610_ (.A1(\fifo_inst.rWrPtrPlus1[3] ),
    .A2(_05867_),
    .B1(_05871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05872_));
 sky130_fd_sc_hd__nor2_1 _12611_ (.A(_05870_),
    .B(_05872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00667_));
 sky130_fd_sc_hd__a21boi_1 _12612_ (.A1(\fifo_inst.rWrPtrPlus1[4] ),
    .A2(_05870_),
    .B1_N(_05860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05873_));
 sky130_fd_sc_hd__o21a_1 _12613_ (.A1(\fifo_inst.rWrPtrPlus1[4] ),
    .A2(_05870_),
    .B1(_05873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00668_));
 sky130_fd_sc_hd__nor2_1 _12614_ (.A(_05279_),
    .B(_05833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05874_));
 sky130_fd_sc_hd__o21a_1 _12615_ (.A1(_05863_),
    .A2(_05874_),
    .B1(_05848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00669_));
 sky130_fd_sc_hd__or2_1 _12616_ (.A(_05865_),
    .B(_05849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05875_));
 sky130_fd_sc_hd__clkbuf_2 _12617_ (.A(_05847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05876_));
 sky130_fd_sc_hd__o211a_1 _12618_ (.A1(_05278_),
    .A2(_05833_),
    .B1(_05875_),
    .C1(_05876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00670_));
 sky130_fd_sc_hd__or2_1 _12619_ (.A(_05342_),
    .B(_05833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05877_));
 sky130_fd_sc_hd__o211a_1 _12620_ (.A1(\fifo_inst.rWrPtrPlus1[2] ),
    .A2(_05849_),
    .B1(_05877_),
    .C1(_05876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00671_));
 sky130_fd_sc_hd__or2_1 _12621_ (.A(_05345_),
    .B(_05832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05878_));
 sky130_fd_sc_hd__o211a_1 _12622_ (.A1(\fifo_inst.rWrPtrPlus1[3] ),
    .A2(_05849_),
    .B1(_05878_),
    .C1(_05876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00672_));
 sky130_fd_sc_hd__or2_1 _12623_ (.A(\fifo_inst.rWrPtr[4] ),
    .B(_05832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05879_));
 sky130_fd_sc_hd__o211a_1 _12624_ (.A1(\fifo_inst.rWrPtrPlus1[4] ),
    .A2(_05849_),
    .B1(_05879_),
    .C1(_05876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00673_));
 sky130_fd_sc_hd__nor2_1 _12625_ (.A(_05842_),
    .B(_05834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05880_));
 sky130_fd_sc_hd__nor2_1 _12626_ (.A(\fifo_inst.rRdPtrPlus1[0] ),
    .B(_04725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05881_));
 sky130_fd_sc_hd__o21ai_1 _12627_ (.A1(_05880_),
    .A2(_05881_),
    .B1(_05848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00674_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12628_ (.A(\fifo_inst.rRdPtrPlus1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05882_));
 sky130_fd_sc_hd__o21ai_1 _12629_ (.A1(_05882_),
    .A2(_05880_),
    .B1(_05847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05883_));
 sky130_fd_sc_hd__a21oi_1 _12630_ (.A1(_05882_),
    .A2(_05880_),
    .B1(_05883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00675_));
 sky130_fd_sc_hd__and3_1 _12631_ (.A(\fifo_inst.rRdPtrPlus1[2] ),
    .B(_05882_),
    .C(_05880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05884_));
 sky130_fd_sc_hd__a31o_1 _12632_ (.A1(_05882_),
    .A2(\fifo_inst.rRdPtrPlus1[0] ),
    .A3(_04724_),
    .B1(\fifo_inst.rRdPtrPlus1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05885_));
 sky130_fd_sc_hd__and3b_1 _12633_ (.A_N(_05884_),
    .B(_05860_),
    .C(_05885_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05886_));
 sky130_fd_sc_hd__clkbuf_1 _12634_ (.A(_05886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00676_));
 sky130_fd_sc_hd__and2_1 _12635_ (.A(\fifo_inst.rRdPtrPlus1[3] ),
    .B(_05884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05887_));
 sky130_fd_sc_hd__o21ai_1 _12636_ (.A1(\fifo_inst.rRdPtrPlus1[3] ),
    .A2(_05884_),
    .B1(_05871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05888_));
 sky130_fd_sc_hd__nor2_1 _12637_ (.A(_05887_),
    .B(_05888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00677_));
 sky130_fd_sc_hd__a21boi_1 _12638_ (.A1(\fifo_inst.rRdPtrPlus1[4] ),
    .A2(_05887_),
    .B1_N(_05860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05889_));
 sky130_fd_sc_hd__o21a_1 _12639_ (.A1(\fifo_inst.rRdPtrPlus1[4] ),
    .A2(_05887_),
    .B1(_05889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00678_));
 sky130_fd_sc_hd__a21o_1 _12640_ (.A1(_04733_),
    .A2(_05834_),
    .B1(_05880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05890_));
 sky130_fd_sc_hd__and2_1 _12641_ (.A(_05847_),
    .B(_05890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05891_));
 sky130_fd_sc_hd__clkbuf_1 _12642_ (.A(_05891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00679_));
 sky130_fd_sc_hd__or2_1 _12643_ (.A(_04737_),
    .B(_04821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05892_));
 sky130_fd_sc_hd__o211a_1 _12644_ (.A1(_05882_),
    .A2(_05835_),
    .B1(_05892_),
    .C1(_05876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00680_));
 sky130_fd_sc_hd__or2_1 _12645_ (.A(_04729_),
    .B(_04821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05893_));
 sky130_fd_sc_hd__o211a_1 _12646_ (.A1(\fifo_inst.rRdPtrPlus1[2] ),
    .A2(_05835_),
    .B1(_05893_),
    .C1(_05871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00681_));
 sky130_fd_sc_hd__or2_1 _12647_ (.A(_05023_),
    .B(_04772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05894_));
 sky130_fd_sc_hd__o211a_1 _12648_ (.A1(\fifo_inst.rRdPtrPlus1[3] ),
    .A2(_05835_),
    .B1(_05894_),
    .C1(_05871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00682_));
 sky130_fd_sc_hd__or2_1 _12649_ (.A(\fifo_inst.rRdPtr[4] ),
    .B(_04772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05895_));
 sky130_fd_sc_hd__o211a_1 _12650_ (.A1(\fifo_inst.rRdPtrPlus1[4] ),
    .A2(_05835_),
    .B1(_05895_),
    .C1(_05871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00683_));
 sky130_fd_sc_hd__dfrtp_1 _12651_ (.CLK(clknet_leaf_19_clk),
    .D(\sa_inst.EOB_Q_o ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12652_ (.CLK(clknet_leaf_20_clk),
    .D(\shift_register[0] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12653_ (.CLK(clknet_leaf_20_clk),
    .D(\shift_register[1] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12654_ (.CLK(clknet_leaf_20_clk),
    .D(\shift_register[2] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12655_ (.CLK(clknet_leaf_20_clk),
    .D(\shift_register[3] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12656_ (.CLK(clknet_leaf_20_clk),
    .D(\shift_register[4] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12657_ (.CLK(clknet_leaf_164_clk),
    .D(\shift_register[5] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12658_ (.CLK(clknet_leaf_164_clk),
    .D(\shift_register[6] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12659_ (.CLK(clknet_leaf_173_clk),
    .D(\shift_register[7] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12660_ (.CLK(clknet_leaf_173_clk),
    .D(\shift_register[8] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12661_ (.CLK(clknet_leaf_173_clk),
    .D(\shift_register[9] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12662_ (.CLK(clknet_leaf_173_clk),
    .D(\shift_register[10] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[11] ));
 sky130_fd_sc_hd__dfxtp_2 _12663_ (.CLK(clknet_leaf_80_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j._12_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._07_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12664_ (.CLK(clknet_leaf_80_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j._12_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._07_[6] ));
 sky130_fd_sc_hd__dfxtp_2 _12665_ (.CLK(clknet_leaf_81_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j._12_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._07_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12666_ (.CLK(clknet_leaf_81_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j._12_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._07_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12667_ (.CLK(clknet_leaf_49_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j._12_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._05_[5] ));
 sky130_fd_sc_hd__dfxtp_2 _12668_ (.CLK(clknet_leaf_53_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j._12_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._05_[6] ));
 sky130_fd_sc_hd__dfxtp_2 _12669_ (.CLK(clknet_leaf_49_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j._12_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._05_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12670_ (.CLK(clknet_leaf_49_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j._12_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._05_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12671_ (.CLK(clknet_leaf_45_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w11_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12672_ (.CLK(clknet_leaf_50_clk),
    .D(_00000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12673_ (.CLK(clknet_leaf_62_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12674_ (.CLK(clknet_leaf_52_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12675_ (.CLK(clknet_leaf_62_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12676_ (.CLK(clknet_leaf_63_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12677_ (.CLK(clknet_leaf_28_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12678_ (.CLK(clknet_leaf_16_clk),
    .D(_00001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._03_ ));
 sky130_fd_sc_hd__dfxtp_1 _12679_ (.CLK(clknet_leaf_120_clk),
    .D(_00002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._03_ ));
 sky130_fd_sc_hd__dfxtp_1 _12680_ (.CLK(clknet_leaf_99_clk),
    .D(_00003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._03_ ));
 sky130_fd_sc_hd__dfxtp_1 _12681_ (.CLK(clknet_leaf_28_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12682_ (.CLK(clknet_leaf_28_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12683_ (.CLK(clknet_leaf_28_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12684_ (.CLK(clknet_leaf_27_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12685_ (.CLK(clknet_leaf_28_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12686_ (.CLK(clknet_leaf_29_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12687_ (.CLK(clknet_leaf_29_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12688_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12689_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12690_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12691_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12692_ (.CLK(clknet_leaf_32_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _12693_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _12694_ (.CLK(clknet_leaf_32_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12695_ (.CLK(clknet_leaf_32_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _12696_ (.CLK(clknet_leaf_32_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _12697_ (.CLK(clknet_leaf_11_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _12698_ (.CLK(clknet_leaf_10_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _12699_ (.CLK(clknet_leaf_11_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _12700_ (.CLK(clknet_leaf_7_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _12701_ (.CLK(clknet_leaf_5_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _12702_ (.CLK(clknet_leaf_5_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _12703_ (.CLK(clknet_leaf_7_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _12704_ (.CLK(clknet_leaf_7_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _12705_ (.CLK(clknet_leaf_7_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _12706_ (.CLK(clknet_leaf_14_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _12707_ (.CLK(clknet_leaf_18_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _12708_ (.CLK(clknet_leaf_26_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[32] ));
 sky130_fd_sc_hd__dfxtp_1 _12709_ (.CLK(clknet_leaf_75_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12710_ (.CLK(clknet_leaf_75_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12711_ (.CLK(clknet_leaf_74_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12712_ (.CLK(clknet_leaf_74_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12713_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12714_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12715_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12716_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12717_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12718_ (.CLK(clknet_leaf_72_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12719_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12720_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12721_ (.CLK(clknet_leaf_108_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12722_ (.CLK(clknet_leaf_111_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12723_ (.CLK(clknet_leaf_111_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12724_ (.CLK(clknet_leaf_111_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12725_ (.CLK(clknet_leaf_111_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _12726_ (.CLK(clknet_leaf_112_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _12727_ (.CLK(clknet_leaf_112_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12728_ (.CLK(clknet_leaf_112_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _12729_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _12730_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _12731_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _12732_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _12733_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _12734_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _12735_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _12736_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _12737_ (.CLK(clknet_leaf_162_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _12738_ (.CLK(clknet_leaf_162_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _12739_ (.CLK(clknet_leaf_162_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _12740_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _12741_ (.CLK(clknet_leaf_70_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[32] ));
 sky130_fd_sc_hd__dfxtp_1 _12742_ (.CLK(clknet_leaf_92_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12743_ (.CLK(clknet_leaf_92_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12744_ (.CLK(clknet_leaf_93_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12745_ (.CLK(clknet_leaf_93_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12746_ (.CLK(clknet_leaf_93_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12747_ (.CLK(clknet_leaf_93_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12748_ (.CLK(clknet_leaf_93_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12749_ (.CLK(clknet_leaf_93_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12750_ (.CLK(clknet_leaf_93_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12751_ (.CLK(clknet_leaf_93_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12752_ (.CLK(clknet_leaf_93_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12753_ (.CLK(clknet_leaf_94_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12754_ (.CLK(clknet_leaf_105_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12755_ (.CLK(clknet_leaf_105_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12756_ (.CLK(clknet_leaf_94_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12757_ (.CLK(clknet_leaf_105_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12758_ (.CLK(clknet_leaf_104_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _12759_ (.CLK(clknet_leaf_104_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _12760_ (.CLK(clknet_leaf_104_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12761_ (.CLK(clknet_leaf_104_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _12762_ (.CLK(clknet_leaf_103_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _12763_ (.CLK(clknet_leaf_103_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _12764_ (.CLK(clknet_leaf_103_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _12765_ (.CLK(clknet_leaf_123_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _12766_ (.CLK(clknet_leaf_123_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _12767_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _12768_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _12769_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _12770_ (.CLK(clknet_leaf_123_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _12771_ (.CLK(clknet_leaf_123_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _12772_ (.CLK(clknet_leaf_123_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _12773_ (.CLK(clknet_leaf_122_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _12774_ (.CLK(clknet_leaf_105_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[32] ));
 sky130_fd_sc_hd__dfxtp_1 _12775_ (.CLK(clknet_leaf_26_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12776_ (.CLK(clknet_leaf_26_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12777_ (.CLK(clknet_leaf_26_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12778_ (.CLK(clknet_leaf_26_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12779_ (.CLK(clknet_leaf_25_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12780_ (.CLK(clknet_leaf_26_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12781_ (.CLK(clknet_leaf_25_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12782_ (.CLK(clknet_leaf_26_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12783_ (.CLK(clknet_leaf_25_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12784_ (.CLK(clknet_leaf_27_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12785_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12786_ (.CLK(clknet_leaf_25_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12787_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12788_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12789_ (.CLK(clknet_leaf_12_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12790_ (.CLK(clknet_leaf_12_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12791_ (.CLK(clknet_leaf_25_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _12792_ (.CLK(clknet_leaf_25_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _12793_ (.CLK(clknet_leaf_25_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12794_ (.CLK(clknet_leaf_13_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _12795_ (.CLK(clknet_leaf_12_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _12796_ (.CLK(clknet_leaf_12_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _12797_ (.CLK(clknet_leaf_12_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _12798_ (.CLK(clknet_leaf_12_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _12799_ (.CLK(clknet_leaf_5_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _12800_ (.CLK(clknet_leaf_5_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _12801_ (.CLK(clknet_leaf_5_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _12802_ (.CLK(clknet_leaf_5_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _12803_ (.CLK(clknet_leaf_5_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _12804_ (.CLK(clknet_leaf_14_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _12805_ (.CLK(clknet_leaf_14_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _12806_ (.CLK(clknet_leaf_19_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _12807_ (.CLK(clknet_leaf_163_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[32] ));
 sky130_fd_sc_hd__dfxtp_1 _12808_ (.CLK(clknet_leaf_116_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12809_ (.CLK(clknet_leaf_117_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12810_ (.CLK(clknet_leaf_116_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12811_ (.CLK(clknet_leaf_117_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12812_ (.CLK(clknet_leaf_116_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12813_ (.CLK(clknet_leaf_117_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12814_ (.CLK(clknet_leaf_117_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12815_ (.CLK(clknet_leaf_118_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12816_ (.CLK(clknet_leaf_118_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12817_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12818_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12819_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12820_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12821_ (.CLK(clknet_leaf_118_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12822_ (.CLK(clknet_leaf_118_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12823_ (.CLK(clknet_leaf_118_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12824_ (.CLK(clknet_leaf_118_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _12825_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _12826_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12827_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _12828_ (.CLK(clknet_leaf_118_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _12829_ (.CLK(clknet_leaf_118_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _12830_ (.CLK(clknet_leaf_118_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _12831_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _12832_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _12833_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _12834_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _12835_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _12836_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _12837_ (.CLK(clknet_leaf_157_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _12838_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _12839_ (.CLK(clknet_leaf_115_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _12840_ (.CLK(clknet_leaf_156_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[32] ));
 sky130_fd_sc_hd__dfxtp_1 _12841_ (.CLK(clknet_leaf_95_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12842_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12843_ (.CLK(clknet_leaf_95_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12844_ (.CLK(clknet_leaf_99_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12845_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12846_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12847_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12848_ (.CLK(clknet_leaf_95_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12849_ (.CLK(clknet_leaf_95_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12850_ (.CLK(clknet_leaf_95_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12851_ (.CLK(clknet_leaf_94_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12852_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12853_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12854_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12855_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12856_ (.CLK(clknet_leaf_102_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12857_ (.CLK(clknet_leaf_101_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _12858_ (.CLK(clknet_leaf_102_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _12859_ (.CLK(clknet_leaf_101_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12860_ (.CLK(clknet_leaf_101_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _12861_ (.CLK(clknet_leaf_101_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _12862_ (.CLK(clknet_leaf_101_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _12863_ (.CLK(clknet_leaf_103_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _12864_ (.CLK(clknet_leaf_103_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _12865_ (.CLK(clknet_leaf_123_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _12866_ (.CLK(clknet_leaf_124_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _12867_ (.CLK(clknet_leaf_124_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _12868_ (.CLK(clknet_leaf_124_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _12869_ (.CLK(clknet_leaf_124_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _12870_ (.CLK(clknet_leaf_124_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _12871_ (.CLK(clknet_leaf_123_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _12872_ (.CLK(clknet_leaf_123_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _12873_ (.CLK(clknet_leaf_131_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.24$func$/openlane/designs/teras/src/pe_s3.v:67$123.$result[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[32] ));
 sky130_fd_sc_hd__dfxtp_1 _12874_ (.CLK(clknet_leaf_79_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._14_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12875_ (.CLK(clknet_leaf_81_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._14_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12876_ (.CLK(clknet_leaf_43_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[0] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12877_ (.CLK(clknet_leaf_42_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[1] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12878_ (.CLK(clknet_leaf_42_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[2] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12879_ (.CLK(clknet_leaf_43_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[3] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12880_ (.CLK(clknet_leaf_43_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[4] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12881_ (.CLK(clknet_leaf_43_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[5] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12882_ (.CLK(clknet_leaf_42_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[6] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12883_ (.CLK(clknet_leaf_37_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[7] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12884_ (.CLK(clknet_leaf_42_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[8] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12885_ (.CLK(clknet_leaf_42_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[9] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12886_ (.CLK(clknet_leaf_37_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[10] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12887_ (.CLK(clknet_leaf_37_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[11] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12888_ (.CLK(clknet_leaf_37_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[12] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12889_ (.CLK(clknet_leaf_35_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[13] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12890_ (.CLK(clknet_leaf_37_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[14] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12891_ (.CLK(clknet_leaf_35_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[15] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12892_ (.CLK(clknet_leaf_35_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[16] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12893_ (.CLK(clknet_leaf_35_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[17] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12894_ (.CLK(clknet_leaf_35_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[18] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12895_ (.CLK(clknet_leaf_35_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[19] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12896_ (.CLK(clknet_leaf_35_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[20] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12897_ (.CLK(clknet_leaf_33_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[21] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12898_ (.CLK(clknet_leaf_34_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[22] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12899_ (.CLK(clknet_leaf_34_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[23] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12900_ (.CLK(clknet_leaf_9_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[24] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12901_ (.CLK(clknet_leaf_9_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[25] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12902_ (.CLK(clknet_leaf_9_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[26] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12903_ (.CLK(clknet_leaf_8_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[27] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12904_ (.CLK(clknet_leaf_8_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[28] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12905_ (.CLK(clknet_leaf_8_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[29] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12906_ (.CLK(clknet_leaf_8_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[30] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12907_ (.CLK(clknet_leaf_9_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._24_[31] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._10_[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12908_ (.CLK(clknet_leaf_36_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._20_ ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._02_ ));
 sky130_fd_sc_hd__dfxtp_4 _12909_ (.CLK(clknet_leaf_47_clk),
    .D(\sa_inst.sak._33_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._10_ ));
 sky130_fd_sc_hd__dfxtp_2 _12910_ (.CLK(clknet_leaf_38_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._17_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._26_ ));
 sky130_fd_sc_hd__dfxtp_1 _12911_ (.CLK(clknet_leaf_35_clk),
    .D(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst._25_ ));
 sky130_fd_sc_hd__dfxtp_1 _12912_ (.CLK(clknet_leaf_167_clk),
    .D(_00004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._02_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12913_ (.CLK(clknet_leaf_173_clk),
    .D(_00005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._02_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12914_ (.CLK(clknet_leaf_161_clk),
    .D(_00006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._02_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12915_ (.CLK(clknet_leaf_160_clk),
    .D(_00007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._02_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12916_ (.CLK(clknet_leaf_160_clk),
    .D(_00008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._02_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12917_ (.CLK(clknet_leaf_159_clk),
    .D(_00009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._02_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12918_ (.CLK(clknet_leaf_159_clk),
    .D(_00010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._02_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12919_ (.CLK(clknet_leaf_41_clk),
    .D(_00011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12920_ (.CLK(clknet_leaf_41_clk),
    .D(_00012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12921_ (.CLK(clknet_leaf_41_clk),
    .D(_00013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12922_ (.CLK(clknet_leaf_41_clk),
    .D(_00014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12923_ (.CLK(clknet_leaf_41_clk),
    .D(_00015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12924_ (.CLK(clknet_leaf_38_clk),
    .D(_00016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12925_ (.CLK(clknet_leaf_38_clk),
    .D(_00017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12926_ (.CLK(clknet_leaf_37_clk),
    .D(_00018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12927_ (.CLK(clknet_leaf_38_clk),
    .D(_00019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12928_ (.CLK(clknet_leaf_38_clk),
    .D(_00020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12929_ (.CLK(clknet_leaf_36_clk),
    .D(_00021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12930_ (.CLK(clknet_leaf_37_clk),
    .D(_00022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12931_ (.CLK(clknet_leaf_36_clk),
    .D(_00023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12932_ (.CLK(clknet_leaf_36_clk),
    .D(_00024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12933_ (.CLK(clknet_leaf_36_clk),
    .D(_00025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12934_ (.CLK(clknet_leaf_36_clk),
    .D(_00026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12935_ (.CLK(clknet_leaf_35_clk),
    .D(_00027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _12936_ (.CLK(clknet_leaf_35_clk),
    .D(_00028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _12937_ (.CLK(clknet_leaf_35_clk),
    .D(_00029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12938_ (.CLK(clknet_leaf_35_clk),
    .D(_00030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _12939_ (.CLK(clknet_leaf_34_clk),
    .D(_00031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _12940_ (.CLK(clknet_leaf_9_clk),
    .D(_00032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _12941_ (.CLK(clknet_leaf_34_clk),
    .D(_00033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _12942_ (.CLK(clknet_leaf_9_clk),
    .D(_00034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _12943_ (.CLK(clknet_leaf_8_clk),
    .D(_00035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _12944_ (.CLK(clknet_leaf_8_clk),
    .D(_00036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _12945_ (.CLK(clknet_leaf_8_clk),
    .D(_00037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _12946_ (.CLK(clknet_leaf_8_clk),
    .D(_00038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _12947_ (.CLK(clknet_leaf_8_clk),
    .D(_00039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _12948_ (.CLK(clknet_leaf_7_clk),
    .D(_00040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _12949_ (.CLK(clknet_leaf_9_clk),
    .D(_00041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _12950_ (.CLK(clknet_leaf_9_clk),
    .D(_00042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _12951_ (.CLK(clknet_leaf_25_clk),
    .D(_00043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[32] ));
 sky130_fd_sc_hd__dfxtp_1 _12952_ (.CLK(clknet_leaf_41_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12953_ (.CLK(clknet_leaf_41_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12954_ (.CLK(clknet_leaf_41_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12955_ (.CLK(clknet_leaf_41_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12956_ (.CLK(clknet_leaf_41_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12957_ (.CLK(clknet_leaf_38_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12958_ (.CLK(clknet_leaf_41_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12959_ (.CLK(clknet_leaf_38_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12960_ (.CLK(clknet_leaf_38_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12961_ (.CLK(clknet_leaf_38_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12962_ (.CLK(clknet_leaf_38_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12963_ (.CLK(clknet_leaf_38_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12964_ (.CLK(clknet_leaf_36_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12965_ (.CLK(clknet_leaf_36_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12966_ (.CLK(clknet_leaf_36_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12967_ (.CLK(clknet_leaf_36_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12968_ (.CLK(clknet_leaf_35_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _12969_ (.CLK(clknet_leaf_33_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _12970_ (.CLK(clknet_leaf_35_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12971_ (.CLK(clknet_leaf_33_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _12972_ (.CLK(clknet_leaf_34_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _12973_ (.CLK(clknet_leaf_34_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _12974_ (.CLK(clknet_leaf_34_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _12975_ (.CLK(clknet_leaf_9_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _12976_ (.CLK(clknet_leaf_8_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _12977_ (.CLK(clknet_leaf_8_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _12978_ (.CLK(clknet_leaf_8_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _12979_ (.CLK(clknet_leaf_8_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _12980_ (.CLK(clknet_leaf_8_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _12981_ (.CLK(clknet_leaf_7_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _12982_ (.CLK(clknet_leaf_9_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _12983_ (.CLK(clknet_leaf_9_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _12984_ (.CLK(clknet_leaf_25_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij._00_[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._40_[32] ));
 sky130_fd_sc_hd__dfxtp_2 _12985_ (.CLK(clknet_leaf_53_clk),
    .D(\sa_inst._05_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._00_[0] ));
 sky130_fd_sc_hd__dfxtp_4 _12986_ (.CLK(clknet_leaf_53_clk),
    .D(\sa_inst._05_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._00_[1] ));
 sky130_fd_sc_hd__dfxtp_2 _12987_ (.CLK(clknet_leaf_61_clk),
    .D(\sa_inst._05_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._00_[2] ));
 sky130_fd_sc_hd__dfxtp_2 _12988_ (.CLK(clknet_leaf_61_clk),
    .D(\sa_inst._05_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._00_[3] ));
 sky130_fd_sc_hd__dfxtp_2 _12989_ (.CLK(clknet_leaf_49_clk),
    .D(\sa_inst._05_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._00_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12990_ (.CLK(clknet_leaf_54_clk),
    .D(\sa_inst._05_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._00_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12991_ (.CLK(clknet_leaf_49_clk),
    .D(\sa_inst._05_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._00_[7] ));
 sky130_fd_sc_hd__dfxtp_2 _12992_ (.CLK(clknet_leaf_49_clk),
    .D(\sa_inst._05_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._00_[8] ));
 sky130_fd_sc_hd__dfxtp_2 _12993_ (.CLK(clknet_leaf_53_clk),
    .D(\sa_inst._05_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._00_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12994_ (.CLK(clknet_leaf_56_clk),
    .D(\sa_inst._05_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._00_[10] ));
 sky130_fd_sc_hd__dfxtp_4 _12995_ (.CLK(clknet_leaf_61_clk),
    .D(\sa_inst._05_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._00_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12996_ (.CLK(clknet_leaf_28_clk),
    .D(\sa_inst._22_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._22_ ));
 sky130_fd_sc_hd__dfxtp_1 _12997_ (.CLK(clknet_leaf_46_clk),
    .D(\sa_inst._01_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._33_ ));
 sky130_fd_sc_hd__dfrtp_1 _12998_ (.CLK(clknet_leaf_52_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[0] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12999_ (.CLK(clknet_leaf_52_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[1] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13000_ (.CLK(clknet_leaf_62_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[2] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13001_ (.CLK(clknet_leaf_62_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[3] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13002_ (.CLK(clknet_leaf_62_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[4] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13003_ (.CLK(clknet_leaf_63_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[5] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13004_ (.CLK(clknet_leaf_63_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[6] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13005_ (.CLK(clknet_leaf_28_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[7] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[7] ));
 sky130_fd_sc_hd__dfrtp_2 _13006_ (.CLK(clknet_leaf_28_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[8] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13007_ (.CLK(clknet_leaf_28_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[9] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[9] ));
 sky130_fd_sc_hd__dfrtp_2 _13008_ (.CLK(clknet_leaf_39_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[10] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13009_ (.CLK(clknet_leaf_29_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[11] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13010_ (.CLK(clknet_leaf_29_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[12] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13011_ (.CLK(clknet_leaf_29_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[13] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13012_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[14] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13013_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[15] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13014_ (.CLK(clknet_leaf_32_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[16] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13015_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[17] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13016_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[18] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13017_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[19] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13018_ (.CLK(clknet_leaf_31_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[20] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13019_ (.CLK(clknet_leaf_12_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[21] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13020_ (.CLK(clknet_leaf_31_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[22] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13021_ (.CLK(clknet_leaf_31_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[23] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[23] ));
 sky130_fd_sc_hd__dfrtp_2 _13022_ (.CLK(clknet_leaf_12_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[24] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[24] ));
 sky130_fd_sc_hd__dfrtp_2 _13023_ (.CLK(clknet_leaf_11_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[25] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13024_ (.CLK(clknet_leaf_11_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[26] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13025_ (.CLK(clknet_leaf_11_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[27] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[27] ));
 sky130_fd_sc_hd__dfrtp_1 _13026_ (.CLK(clknet_leaf_14_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[28] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[28] ));
 sky130_fd_sc_hd__dfrtp_1 _13027_ (.CLK(clknet_leaf_11_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[29] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[29] ));
 sky130_fd_sc_hd__dfrtp_1 _13028_ (.CLK(clknet_leaf_5_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[30] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[30] ));
 sky130_fd_sc_hd__dfrtp_1 _13029_ (.CLK(clknet_leaf_14_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._24_[31] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._10_[31] ));
 sky130_fd_sc_hd__dfrtp_1 _13030_ (.CLK(clknet_leaf_27_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._20_ ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._02_ ));
 sky130_fd_sc_hd__dfxtp_1 _13031_ (.CLK(clknet_leaf_31_clk),
    .D(\sa_inst.sak._10_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._05_ ));
 sky130_fd_sc_hd__dfxtp_1 _13032_ (.CLK(clknet_leaf_27_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._17_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._26_ ));
 sky130_fd_sc_hd__dfxtp_1 _13033_ (.CLK(clknet_leaf_27_clk),
    .D(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._25_ ));
 sky130_fd_sc_hd__dfxtp_1 _13034_ (.CLK(clknet_leaf_41_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._08_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._22_ ));
 sky130_fd_sc_hd__dfxtp_1 _13035_ (.CLK(clknet_leaf_27_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._02_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._11_ ));
 sky130_fd_sc_hd__dfxtp_1 _13036_ (.CLK(clknet_leaf_50_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._01_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._00_ ));
 sky130_fd_sc_hd__dfxtp_1 _13037_ (.CLK(clknet_leaf_50_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._08_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13038_ (.CLK(clknet_leaf_41_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._08_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13039_ (.CLK(clknet_leaf_41_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst._08_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13040_ (.CLK(clknet_leaf_61_clk),
    .D(_00044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13041_ (.CLK(clknet_leaf_61_clk),
    .D(_00045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13042_ (.CLK(clknet_leaf_62_clk),
    .D(_00046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13043_ (.CLK(clknet_leaf_62_clk),
    .D(_00047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13044_ (.CLK(clknet_leaf_64_clk),
    .D(_00048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13045_ (.CLK(clknet_leaf_64_clk),
    .D(_00049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13046_ (.CLK(clknet_leaf_64_clk),
    .D(_00050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13047_ (.CLK(clknet_leaf_64_clk),
    .D(_00051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13048_ (.CLK(clknet_leaf_64_clk),
    .D(_00052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13049_ (.CLK(clknet_leaf_64_clk),
    .D(_00053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13050_ (.CLK(clknet_leaf_64_clk),
    .D(_00054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13051_ (.CLK(clknet_leaf_27_clk),
    .D(_00055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13052_ (.CLK(clknet_leaf_26_clk),
    .D(_00056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13053_ (.CLK(clknet_leaf_26_clk),
    .D(_00057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13054_ (.CLK(clknet_leaf_26_clk),
    .D(_00058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13055_ (.CLK(clknet_leaf_26_clk),
    .D(_00059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13056_ (.CLK(clknet_leaf_24_clk),
    .D(_00060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13057_ (.CLK(clknet_leaf_24_clk),
    .D(_00061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13058_ (.CLK(clknet_leaf_24_clk),
    .D(_00062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13059_ (.CLK(clknet_leaf_24_clk),
    .D(_00063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13060_ (.CLK(clknet_leaf_19_clk),
    .D(_00064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13061_ (.CLK(clknet_leaf_19_clk),
    .D(_00065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13062_ (.CLK(clknet_leaf_19_clk),
    .D(_00066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13063_ (.CLK(clknet_leaf_19_clk),
    .D(_00067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13064_ (.CLK(clknet_leaf_20_clk),
    .D(_00068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13065_ (.CLK(clknet_leaf_20_clk),
    .D(_00069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13066_ (.CLK(clknet_leaf_20_clk),
    .D(_00070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13067_ (.CLK(clknet_leaf_164_clk),
    .D(_00071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13068_ (.CLK(clknet_leaf_164_clk),
    .D(_00072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13069_ (.CLK(clknet_leaf_20_clk),
    .D(_00073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13070_ (.CLK(clknet_leaf_20_clk),
    .D(_00074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13071_ (.CLK(clknet_leaf_164_clk),
    .D(_00075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13072_ (.CLK(clknet_leaf_27_clk),
    .D(_00076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[32] ));
 sky130_fd_sc_hd__dfxtp_1 _13073_ (.CLK(clknet_leaf_60_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13074_ (.CLK(clknet_leaf_61_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13075_ (.CLK(clknet_leaf_59_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13076_ (.CLK(clknet_leaf_59_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13077_ (.CLK(clknet_leaf_64_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13078_ (.CLK(clknet_leaf_64_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13079_ (.CLK(clknet_leaf_71_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13080_ (.CLK(clknet_leaf_71_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13081_ (.CLK(clknet_leaf_71_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13082_ (.CLK(clknet_leaf_64_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13083_ (.CLK(clknet_leaf_64_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13084_ (.CLK(clknet_leaf_64_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13085_ (.CLK(clknet_leaf_26_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13086_ (.CLK(clknet_leaf_26_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13087_ (.CLK(clknet_leaf_70_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13088_ (.CLK(clknet_leaf_23_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13089_ (.CLK(clknet_leaf_23_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13090_ (.CLK(clknet_leaf_24_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13091_ (.CLK(clknet_leaf_24_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13092_ (.CLK(clknet_leaf_24_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13093_ (.CLK(clknet_leaf_19_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13094_ (.CLK(clknet_leaf_19_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13095_ (.CLK(clknet_leaf_19_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13096_ (.CLK(clknet_leaf_19_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13097_ (.CLK(clknet_leaf_164_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13098_ (.CLK(clknet_leaf_20_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13099_ (.CLK(clknet_leaf_20_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13100_ (.CLK(clknet_leaf_164_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13101_ (.CLK(clknet_leaf_164_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13102_ (.CLK(clknet_leaf_164_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13103_ (.CLK(clknet_leaf_164_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13104_ (.CLK(clknet_leaf_163_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13105_ (.CLK(clknet_leaf_27_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij._00_[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._01_[32] ));
 sky130_fd_sc_hd__dfxtp_2 _13106_ (.CLK(clknet_leaf_53_clk),
    .D(\sa_inst.sak._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._08_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13107_ (.CLK(clknet_leaf_53_clk),
    .D(\sa_inst.sak._00_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._08_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13108_ (.CLK(clknet_leaf_61_clk),
    .D(\sa_inst.sak._00_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._08_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13109_ (.CLK(clknet_leaf_61_clk),
    .D(\sa_inst.sak._00_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._08_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13110_ (.CLK(clknet_leaf_56_clk),
    .D(\sa_inst.sak._00_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._08_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13111_ (.CLK(clknet_leaf_57_clk),
    .D(\sa_inst.sak._00_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._08_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13112_ (.CLK(clknet_leaf_57_clk),
    .D(\sa_inst.sak._00_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._08_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13113_ (.CLK(clknet_leaf_56_clk),
    .D(\sa_inst.sak._00_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._08_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13114_ (.CLK(clknet_leaf_56_clk),
    .D(\sa_inst.sak._00_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._08_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13115_ (.CLK(clknet_leaf_56_clk),
    .D(\sa_inst.sak._00_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._08_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13116_ (.CLK(clknet_leaf_58_clk),
    .D(\sa_inst.sak._00_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._08_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13117_ (.CLK(clknet_leaf_67_clk),
    .D(\sa_inst.sak._00_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._08_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13118_ (.CLK(clknet_leaf_78_clk),
    .D(\sa_inst._06_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._07_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13119_ (.CLK(clknet_leaf_60_clk),
    .D(\sa_inst._06_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._07_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13120_ (.CLK(clknet_leaf_77_clk),
    .D(\sa_inst._06_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._07_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13121_ (.CLK(clknet_leaf_77_clk),
    .D(\sa_inst._06_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._07_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13122_ (.CLK(clknet_leaf_58_clk),
    .D(\sa_inst._06_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._07_[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13123_ (.CLK(clknet_leaf_56_clk),
    .D(\sa_inst._06_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._07_[5] ));
 sky130_fd_sc_hd__dfxtp_2 _13124_ (.CLK(clknet_leaf_56_clk),
    .D(\sa_inst._06_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._07_[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13125_ (.CLK(clknet_leaf_56_clk),
    .D(\sa_inst._06_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._07_[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13126_ (.CLK(clknet_leaf_56_clk),
    .D(\sa_inst._06_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._07_[8] ));
 sky130_fd_sc_hd__dfxtp_2 _13127_ (.CLK(clknet_leaf_56_clk),
    .D(\sa_inst._06_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._07_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13128_ (.CLK(clknet_leaf_83_clk),
    .D(\sa_inst._06_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._07_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13129_ (.CLK(clknet_leaf_71_clk),
    .D(\sa_inst._06_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._07_[11] ));
 sky130_fd_sc_hd__dfxtp_2 _13130_ (.CLK(clknet_leaf_27_clk),
    .D(\sa_inst.sak._22_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._09_ ));
 sky130_fd_sc_hd__dfrtp_1 _13131_ (.CLK(clknet_leaf_60_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[0] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13132_ (.CLK(clknet_leaf_60_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[1] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13133_ (.CLK(clknet_leaf_60_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[2] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13134_ (.CLK(clknet_leaf_65_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[3] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13135_ (.CLK(clknet_leaf_65_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[4] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13136_ (.CLK(clknet_leaf_66_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[5] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13137_ (.CLK(clknet_leaf_66_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[6] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13138_ (.CLK(clknet_leaf_71_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[7] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13139_ (.CLK(clknet_leaf_71_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[8] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13140_ (.CLK(clknet_leaf_67_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[9] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13141_ (.CLK(clknet_leaf_67_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[10] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13142_ (.CLK(clknet_leaf_67_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[11] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13143_ (.CLK(clknet_leaf_68_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[12] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13144_ (.CLK(clknet_leaf_68_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[13] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[13] ));
 sky130_fd_sc_hd__dfrtp_2 _13145_ (.CLK(clknet_leaf_68_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[14] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13146_ (.CLK(clknet_leaf_68_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[15] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13147_ (.CLK(clknet_leaf_69_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[16] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13148_ (.CLK(clknet_leaf_68_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[17] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13149_ (.CLK(clknet_leaf_69_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[18] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13150_ (.CLK(clknet_leaf_69_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[19] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13151_ (.CLK(clknet_leaf_69_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[20] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13152_ (.CLK(clknet_leaf_112_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[21] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13153_ (.CLK(clknet_leaf_21_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[22] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13154_ (.CLK(clknet_leaf_113_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[23] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[23] ));
 sky130_fd_sc_hd__dfrtp_2 _13155_ (.CLK(clknet_leaf_163_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[24] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13156_ (.CLK(clknet_leaf_163_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[25] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13157_ (.CLK(clknet_leaf_21_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[26] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13158_ (.CLK(clknet_leaf_163_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[27] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[27] ));
 sky130_fd_sc_hd__dfrtp_1 _13159_ (.CLK(clknet_leaf_21_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[28] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[28] ));
 sky130_fd_sc_hd__dfrtp_1 _13160_ (.CLK(clknet_leaf_22_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[29] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[29] ));
 sky130_fd_sc_hd__dfrtp_1 _13161_ (.CLK(clknet_leaf_22_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[30] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[30] ));
 sky130_fd_sc_hd__dfrtp_1 _13162_ (.CLK(clknet_leaf_22_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._24_[31] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._10_[31] ));
 sky130_fd_sc_hd__dfrtp_1 _13163_ (.CLK(clknet_leaf_70_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._20_ ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._02_ ));
 sky130_fd_sc_hd__dfxtp_1 _13164_ (.CLK(clknet_leaf_24_clk),
    .D(\sa_inst.sak._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._21_ ));
 sky130_fd_sc_hd__dfxtp_1 _13165_ (.CLK(clknet_leaf_70_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._17_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._26_ ));
 sky130_fd_sc_hd__dfxtp_1 _13166_ (.CLK(clknet_leaf_68_clk),
    .D(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._25_ ));
 sky130_fd_sc_hd__dfxtp_1 _13167_ (.CLK(clknet_leaf_60_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._08_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._22_ ));
 sky130_fd_sc_hd__dfxtp_1 _13168_ (.CLK(clknet_leaf_70_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._02_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._11_ ));
 sky130_fd_sc_hd__dfxtp_1 _13169_ (.CLK(clknet_leaf_58_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._01_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._00_ ));
 sky130_fd_sc_hd__dfxtp_1 _13170_ (.CLK(clknet_leaf_58_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._08_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ));
 sky130_fd_sc_hd__dfxtp_2 _13171_ (.CLK(clknet_leaf_58_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._08_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13172_ (.CLK(clknet_leaf_60_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst._08_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13173_ (.CLK(clknet_leaf_75_clk),
    .D(_00077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13174_ (.CLK(clknet_leaf_75_clk),
    .D(_00078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13175_ (.CLK(clknet_leaf_76_clk),
    .D(_00079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13176_ (.CLK(clknet_leaf_76_clk),
    .D(_00080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13177_ (.CLK(clknet_leaf_73_clk),
    .D(_00081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13178_ (.CLK(clknet_leaf_73_clk),
    .D(_00082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13179_ (.CLK(clknet_leaf_73_clk),
    .D(_00083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13180_ (.CLK(clknet_leaf_73_clk),
    .D(_00084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13181_ (.CLK(clknet_leaf_71_clk),
    .D(_00085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13182_ (.CLK(clknet_leaf_70_clk),
    .D(_00086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13183_ (.CLK(clknet_leaf_70_clk),
    .D(_00087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13184_ (.CLK(clknet_leaf_70_clk),
    .D(_00088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13185_ (.CLK(clknet_leaf_70_clk),
    .D(_00089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13186_ (.CLK(clknet_leaf_70_clk),
    .D(_00090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13187_ (.CLK(clknet_leaf_70_clk),
    .D(_00091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13188_ (.CLK(clknet_leaf_70_clk),
    .D(_00092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13189_ (.CLK(clknet_leaf_111_clk),
    .D(_00093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13190_ (.CLK(clknet_leaf_70_clk),
    .D(_00094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13191_ (.CLK(clknet_leaf_111_clk),
    .D(_00095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13192_ (.CLK(clknet_leaf_111_clk),
    .D(_00096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13193_ (.CLK(clknet_leaf_109_clk),
    .D(_00097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13194_ (.CLK(clknet_leaf_111_clk),
    .D(_00098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13195_ (.CLK(clknet_leaf_111_clk),
    .D(_00099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13196_ (.CLK(clknet_leaf_112_clk),
    .D(_00100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13197_ (.CLK(clknet_leaf_114_clk),
    .D(_00101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13198_ (.CLK(clknet_leaf_114_clk),
    .D(_00102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13199_ (.CLK(clknet_leaf_162_clk),
    .D(_00103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13200_ (.CLK(clknet_leaf_114_clk),
    .D(_00104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13201_ (.CLK(clknet_leaf_114_clk),
    .D(_00105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13202_ (.CLK(clknet_leaf_112_clk),
    .D(_00106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13203_ (.CLK(clknet_leaf_112_clk),
    .D(_00107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13204_ (.CLK(clknet_leaf_111_clk),
    .D(_00108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13205_ (.CLK(clknet_leaf_108_clk),
    .D(_00109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[32] ));
 sky130_fd_sc_hd__dfxtp_1 _13206_ (.CLK(clknet_leaf_75_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13207_ (.CLK(clknet_leaf_75_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13208_ (.CLK(clknet_leaf_74_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13209_ (.CLK(clknet_leaf_74_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13210_ (.CLK(clknet_leaf_74_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13211_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13212_ (.CLK(clknet_leaf_93_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13213_ (.CLK(clknet_leaf_106_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13214_ (.CLK(clknet_leaf_71_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13215_ (.CLK(clknet_leaf_72_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13216_ (.CLK(clknet_leaf_70_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13217_ (.CLK(clknet_leaf_107_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13218_ (.CLK(clknet_leaf_70_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13219_ (.CLK(clknet_leaf_70_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13220_ (.CLK(clknet_leaf_111_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13221_ (.CLK(clknet_leaf_70_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13222_ (.CLK(clknet_leaf_111_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13223_ (.CLK(clknet_leaf_111_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13224_ (.CLK(clknet_leaf_111_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13225_ (.CLK(clknet_leaf_109_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13226_ (.CLK(clknet_leaf_109_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13227_ (.CLK(clknet_leaf_109_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13228_ (.CLK(clknet_leaf_109_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13229_ (.CLK(clknet_leaf_110_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13230_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13231_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13232_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13233_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13234_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13235_ (.CLK(clknet_leaf_111_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13236_ (.CLK(clknet_leaf_109_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13237_ (.CLK(clknet_leaf_109_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13238_ (.CLK(clknet_leaf_107_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij._00_[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._06_[32] ));
 sky130_fd_sc_hd__dfxtp_2 _13239_ (.CLK(clknet_leaf_84_clk),
    .D(\sa_inst._07_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._03_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13240_ (.CLK(clknet_leaf_84_clk),
    .D(\sa_inst._07_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._03_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13241_ (.CLK(clknet_leaf_84_clk),
    .D(\sa_inst._07_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._03_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13242_ (.CLK(clknet_leaf_84_clk),
    .D(\sa_inst._07_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._03_[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13243_ (.CLK(clknet_leaf_80_clk),
    .D(\sa_inst._07_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._03_[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13244_ (.CLK(clknet_leaf_82_clk),
    .D(\sa_inst._07_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._03_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13245_ (.CLK(clknet_leaf_81_clk),
    .D(\sa_inst._07_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._03_[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13246_ (.CLK(clknet_leaf_82_clk),
    .D(\sa_inst._07_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._03_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13247_ (.CLK(clknet_leaf_82_clk),
    .D(\sa_inst._07_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._03_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13248_ (.CLK(clknet_leaf_82_clk),
    .D(\sa_inst._07_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._03_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13249_ (.CLK(clknet_leaf_83_clk),
    .D(\sa_inst._07_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._03_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13250_ (.CLK(clknet_leaf_72_clk),
    .D(\sa_inst._07_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._03_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13251_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak._09_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._04_ ));
 sky130_fd_sc_hd__dfrtp_1 _13252_ (.CLK(clknet_leaf_51_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[0] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13253_ (.CLK(clknet_leaf_51_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[1] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13254_ (.CLK(clknet_leaf_40_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[2] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13255_ (.CLK(clknet_leaf_40_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[3] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13256_ (.CLK(clknet_leaf_63_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[4] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[4] ));
 sky130_fd_sc_hd__dfrtp_2 _13257_ (.CLK(clknet_leaf_28_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[5] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[5] ));
 sky130_fd_sc_hd__dfrtp_4 _13258_ (.CLK(clknet_leaf_40_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[6] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13259_ (.CLK(clknet_leaf_39_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[7] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13260_ (.CLK(clknet_leaf_39_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[8] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13261_ (.CLK(clknet_leaf_38_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[9] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13262_ (.CLK(clknet_leaf_38_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[10] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13263_ (.CLK(clknet_leaf_38_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[11] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13264_ (.CLK(clknet_leaf_39_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[12] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13265_ (.CLK(clknet_leaf_36_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[13] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13266_ (.CLK(clknet_leaf_32_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[14] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13267_ (.CLK(clknet_leaf_33_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[15] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13268_ (.CLK(clknet_leaf_33_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[16] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13269_ (.CLK(clknet_leaf_33_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[17] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13270_ (.CLK(clknet_leaf_33_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[18] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13271_ (.CLK(clknet_leaf_33_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[19] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13272_ (.CLK(clknet_leaf_33_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[20] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13273_ (.CLK(clknet_leaf_33_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[21] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13274_ (.CLK(clknet_leaf_9_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[22] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13275_ (.CLK(clknet_leaf_10_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[23] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[23] ));
 sky130_fd_sc_hd__dfrtp_2 _13276_ (.CLK(clknet_leaf_10_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[24] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[24] ));
 sky130_fd_sc_hd__dfrtp_2 _13277_ (.CLK(clknet_leaf_10_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[25] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13278_ (.CLK(clknet_leaf_8_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[26] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13279_ (.CLK(clknet_leaf_7_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[27] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[27] ));
 sky130_fd_sc_hd__dfrtp_1 _13280_ (.CLK(clknet_leaf_8_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[28] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[28] ));
 sky130_fd_sc_hd__dfrtp_1 _13281_ (.CLK(clknet_leaf_7_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[29] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[29] ));
 sky130_fd_sc_hd__dfrtp_1 _13282_ (.CLK(clknet_leaf_7_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[30] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[30] ));
 sky130_fd_sc_hd__dfrtp_1 _13283_ (.CLK(clknet_leaf_10_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._24_[31] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._10_[31] ));
 sky130_fd_sc_hd__dfrtp_1 _13284_ (.CLK(clknet_leaf_27_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij.s3fdp_inst._20_ ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:1.pe_ij._02_ ));
 sky130_fd_sc_hd__dfxtp_1 _13285_ (.CLK(clknet_leaf_62_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13286_ (.CLK(clknet_leaf_62_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13287_ (.CLK(clknet_leaf_62_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13288_ (.CLK(clknet_leaf_62_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13289_ (.CLK(clknet_leaf_28_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13290_ (.CLK(clknet_leaf_28_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13291_ (.CLK(clknet_leaf_28_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13292_ (.CLK(clknet_leaf_28_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13293_ (.CLK(clknet_leaf_27_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13294_ (.CLK(clknet_leaf_27_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13295_ (.CLK(clknet_leaf_29_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13296_ (.CLK(clknet_leaf_28_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13297_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13298_ (.CLK(clknet_leaf_29_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13299_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13300_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13301_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13302_ (.CLK(clknet_leaf_25_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13303_ (.CLK(clknet_leaf_30_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13304_ (.CLK(clknet_leaf_32_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13305_ (.CLK(clknet_leaf_12_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13306_ (.CLK(clknet_leaf_12_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13307_ (.CLK(clknet_leaf_12_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13308_ (.CLK(clknet_leaf_12_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13309_ (.CLK(clknet_leaf_5_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13310_ (.CLK(clknet_leaf_5_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13311_ (.CLK(clknet_leaf_5_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13312_ (.CLK(clknet_leaf_5_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13313_ (.CLK(clknet_leaf_5_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13314_ (.CLK(clknet_leaf_7_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13315_ (.CLK(clknet_leaf_14_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13316_ (.CLK(clknet_leaf_18_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13317_ (.CLK(clknet_leaf_26_clk),
    .D(\sa_inst.sak.rows:2.cols:1.pe_ij._00_[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._12_[32] ));
 sky130_fd_sc_hd__dfxtp_4 _13318_ (.CLK(clknet_leaf_183_clk),
    .D(_00110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_4 _13319_ (.CLK(clknet_leaf_183_clk),
    .D(_00111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_2 _13320_ (.CLK(clknet_leaf_183_clk),
    .D(_00112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _13321_ (.CLK(clknet_leaf_183_clk),
    .D(_00113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_4 _13322_ (.CLK(clknet_leaf_183_clk),
    .D(_00114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_4 _13323_ (.CLK(clknet_leaf_155_clk),
    .D(_00115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _13324_ (.CLK(clknet_leaf_154_clk),
    .D(_00116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_4 _13325_ (.CLK(clknet_leaf_156_clk),
    .D(_00117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_4 _13326_ (.CLK(clknet_leaf_156_clk),
    .D(_00118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_4 _13327_ (.CLK(clknet_leaf_154_clk),
    .D(_00119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_4 _13328_ (.CLK(clknet_leaf_152_clk),
    .D(_00120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_4 _13329_ (.CLK(clknet_leaf_152_clk),
    .D(_00121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_2 _13330_ (.CLK(clknet_leaf_145_clk),
    .D(_00122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_1 _13331_ (.CLK(clknet_leaf_148_clk),
    .D(_00123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_4 _13332_ (.CLK(clknet_leaf_144_clk),
    .D(_00124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_4 _13333_ (.CLK(clknet_leaf_185_clk),
    .D(_00125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_4 _13334_ (.CLK(clknet_leaf_185_clk),
    .D(_00126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_4 _13335_ (.CLK(clknet_leaf_1_clk),
    .D(_00127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_2 _13336_ (.CLK(clknet_leaf_1_clk),
    .D(_00128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_4 _13337_ (.CLK(clknet_leaf_1_clk),
    .D(_00129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_2 _13338_ (.CLK(clknet_leaf_192_clk),
    .D(_00130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_1 _13339_ (.CLK(clknet_leaf_192_clk),
    .D(_00131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_4 _13340_ (.CLK(clknet_leaf_186_clk),
    .D(_00132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_1 _13341_ (.CLK(clknet_leaf_186_clk),
    .D(_00133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _13342_ (.CLK(clknet_leaf_47_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13343_ (.CLK(clknet_leaf_47_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13344_ (.CLK(clknet_leaf_47_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13345_ (.CLK(clknet_leaf_47_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13346_ (.CLK(clknet_leaf_47_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13347_ (.CLK(clknet_leaf_48_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13348_ (.CLK(clknet_leaf_47_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13349_ (.CLK(clknet_leaf_47_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13350_ (.CLK(clknet_leaf_50_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13351_ (.CLK(clknet_leaf_49_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13352_ (.CLK(clknet_leaf_50_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13353_ (.CLK(clknet_leaf_50_clk),
    .D(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13354_ (.CLK(clknet_leaf_77_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[0] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13355_ (.CLK(clknet_leaf_77_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[1] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13356_ (.CLK(clknet_leaf_76_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[2] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13357_ (.CLK(clknet_leaf_77_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[3] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13358_ (.CLK(clknet_leaf_71_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[4] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13359_ (.CLK(clknet_leaf_66_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[5] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13360_ (.CLK(clknet_leaf_71_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[6] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13361_ (.CLK(clknet_leaf_71_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[7] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13362_ (.CLK(clknet_leaf_76_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[8] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13363_ (.CLK(clknet_leaf_72_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[9] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13364_ (.CLK(clknet_leaf_72_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[10] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13365_ (.CLK(clknet_leaf_72_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[11] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13366_ (.CLK(clknet_leaf_72_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[12] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13367_ (.CLK(clknet_leaf_70_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[13] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13368_ (.CLK(clknet_leaf_70_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[14] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13369_ (.CLK(clknet_leaf_107_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[15] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13370_ (.CLK(clknet_leaf_69_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[16] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13371_ (.CLK(clknet_leaf_112_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[17] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13372_ (.CLK(clknet_leaf_112_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[18] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13373_ (.CLK(clknet_leaf_113_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[19] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13374_ (.CLK(clknet_leaf_113_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[20] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13375_ (.CLK(clknet_leaf_113_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[21] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13376_ (.CLK(clknet_leaf_163_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[22] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13377_ (.CLK(clknet_leaf_113_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[23] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13378_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[24] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13379_ (.CLK(clknet_leaf_162_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[25] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13380_ (.CLK(clknet_leaf_162_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[26] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13381_ (.CLK(clknet_leaf_162_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[27] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[27] ));
 sky130_fd_sc_hd__dfrtp_1 _13382_ (.CLK(clknet_leaf_163_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[28] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[28] ));
 sky130_fd_sc_hd__dfrtp_1 _13383_ (.CLK(clknet_leaf_162_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[29] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[29] ));
 sky130_fd_sc_hd__dfrtp_1 _13384_ (.CLK(clknet_leaf_163_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[30] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[30] ));
 sky130_fd_sc_hd__dfrtp_1 _13385_ (.CLK(clknet_leaf_163_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._24_[31] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._10_[31] ));
 sky130_fd_sc_hd__dfrtp_1 _13386_ (.CLK(clknet_leaf_70_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._20_ ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij._02_ ));
 sky130_fd_sc_hd__dfxtp_1 _13387_ (.CLK(clknet_leaf_70_clk),
    .D(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst._25_ ));
 sky130_fd_sc_hd__dfxtp_1 _13388_ (.CLK(clknet_leaf_52_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._14_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13389_ (.CLK(clknet_leaf_51_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._14_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13390_ (.CLK(clknet_leaf_77_clk),
    .D(_00134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13391_ (.CLK(clknet_leaf_75_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13392_ (.CLK(clknet_leaf_75_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13393_ (.CLK(clknet_leaf_74_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13394_ (.CLK(clknet_leaf_74_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13395_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13396_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13397_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13398_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13399_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13400_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13401_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13402_ (.CLK(clknet_leaf_107_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13403_ (.CLK(clknet_leaf_108_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13404_ (.CLK(clknet_leaf_111_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13405_ (.CLK(clknet_leaf_108_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13406_ (.CLK(clknet_leaf_108_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13407_ (.CLK(clknet_leaf_111_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13408_ (.CLK(clknet_leaf_111_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13409_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13410_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13411_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13412_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13413_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13414_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13415_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13416_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13417_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13418_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13419_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13420_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13421_ (.CLK(clknet_leaf_162_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13422_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13423_ (.CLK(clknet_leaf_70_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij._00_[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._17_[32] ));
 sky130_fd_sc_hd__dfxtp_1 _13424_ (.CLK(clknet_leaf_78_clk),
    .D(\sa_inst.sak._07_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._13_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13425_ (.CLK(clknet_leaf_78_clk),
    .D(\sa_inst.sak._07_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._13_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13426_ (.CLK(clknet_leaf_77_clk),
    .D(\sa_inst.sak._07_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._13_[2] ));
 sky130_fd_sc_hd__dfxtp_2 _13427_ (.CLK(clknet_leaf_78_clk),
    .D(\sa_inst.sak._07_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._13_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13428_ (.CLK(clknet_leaf_82_clk),
    .D(\sa_inst.sak._07_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._13_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13429_ (.CLK(clknet_leaf_83_clk),
    .D(\sa_inst.sak._07_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._13_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13430_ (.CLK(clknet_leaf_83_clk),
    .D(\sa_inst.sak._07_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._13_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13431_ (.CLK(clknet_leaf_83_clk),
    .D(\sa_inst.sak._07_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._13_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13432_ (.CLK(clknet_leaf_83_clk),
    .D(\sa_inst.sak._07_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._13_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13433_ (.CLK(clknet_leaf_83_clk),
    .D(\sa_inst.sak._07_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._13_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13434_ (.CLK(clknet_leaf_71_clk),
    .D(\sa_inst.sak._07_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._13_[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13435_ (.CLK(clknet_leaf_85_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[0] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13436_ (.CLK(clknet_leaf_84_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[1] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13437_ (.CLK(clknet_leaf_74_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[2] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13438_ (.CLK(clknet_leaf_85_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[3] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13439_ (.CLK(clknet_leaf_106_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[4] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13440_ (.CLK(clknet_leaf_93_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[5] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13441_ (.CLK(clknet_leaf_93_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[6] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13442_ (.CLK(clknet_leaf_106_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[7] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13443_ (.CLK(clknet_leaf_93_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[8] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13444_ (.CLK(clknet_leaf_93_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[9] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13445_ (.CLK(clknet_leaf_106_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[10] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13446_ (.CLK(clknet_leaf_106_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[11] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13447_ (.CLK(clknet_leaf_105_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[12] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13448_ (.CLK(clknet_leaf_104_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[13] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13449_ (.CLK(clknet_leaf_105_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[14] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13450_ (.CLK(clknet_leaf_104_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[15] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13451_ (.CLK(clknet_leaf_103_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[16] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13452_ (.CLK(clknet_leaf_104_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[17] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13453_ (.CLK(clknet_leaf_109_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[18] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13454_ (.CLK(clknet_leaf_109_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[19] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13455_ (.CLK(clknet_leaf_103_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[20] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13456_ (.CLK(clknet_leaf_109_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[21] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13457_ (.CLK(clknet_leaf_109_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[22] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13458_ (.CLK(clknet_leaf_122_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[23] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[23] ));
 sky130_fd_sc_hd__dfrtp_2 _13459_ (.CLK(clknet_leaf_122_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[24] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[24] ));
 sky130_fd_sc_hd__dfrtp_2 _13460_ (.CLK(clknet_leaf_123_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[25] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13461_ (.CLK(clknet_leaf_122_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[26] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13462_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[27] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[27] ));
 sky130_fd_sc_hd__dfrtp_1 _13463_ (.CLK(clknet_leaf_116_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[28] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[28] ));
 sky130_fd_sc_hd__dfrtp_1 _13464_ (.CLK(clknet_leaf_116_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[29] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[29] ));
 sky130_fd_sc_hd__dfrtp_1 _13465_ (.CLK(clknet_leaf_116_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[30] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[30] ));
 sky130_fd_sc_hd__dfrtp_1 _13466_ (.CLK(clknet_leaf_116_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._24_[31] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._10_[31] ));
 sky130_fd_sc_hd__dfrtp_1 _13467_ (.CLK(clknet_leaf_107_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._20_ ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij._02_ ));
 sky130_fd_sc_hd__dfxtp_4 _13468_ (.CLK(clknet_leaf_24_clk),
    .D(\sa_inst.sak._21_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.EOB_Q_o ));
 sky130_fd_sc_hd__dfxtp_1 _13469_ (.CLK(clknet_leaf_107_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._17_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._26_ ));
 sky130_fd_sc_hd__dfxtp_1 _13470_ (.CLK(clknet_leaf_107_clk),
    .D(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._25_ ));
 sky130_fd_sc_hd__dfxtp_1 _13471_ (.CLK(clknet_leaf_85_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._08_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._22_ ));
 sky130_fd_sc_hd__dfxtp_1 _13472_ (.CLK(clknet_leaf_107_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._02_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._11_ ));
 sky130_fd_sc_hd__dfxtp_1 _13473_ (.CLK(clknet_leaf_86_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._01_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._00_ ));
 sky130_fd_sc_hd__dfxtp_1 _13474_ (.CLK(clknet_leaf_85_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._08_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ));
 sky130_fd_sc_hd__dfxtp_2 _13475_ (.CLK(clknet_leaf_85_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._08_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13476_ (.CLK(clknet_leaf_85_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst._08_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13477_ (.CLK(clknet_leaf_75_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w11_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13478_ (.CLK(clknet_leaf_92_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13479_ (.CLK(clknet_leaf_91_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13480_ (.CLK(clknet_leaf_91_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13481_ (.CLK(clknet_leaf_92_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13482_ (.CLK(clknet_leaf_93_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13483_ (.CLK(clknet_leaf_91_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13484_ (.CLK(clknet_leaf_95_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13485_ (.CLK(clknet_leaf_95_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13486_ (.CLK(clknet_leaf_95_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13487_ (.CLK(clknet_leaf_95_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13488_ (.CLK(clknet_leaf_94_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13489_ (.CLK(clknet_leaf_94_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13490_ (.CLK(clknet_leaf_94_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13491_ (.CLK(clknet_leaf_94_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13492_ (.CLK(clknet_leaf_94_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13493_ (.CLK(clknet_leaf_105_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13494_ (.CLK(clknet_leaf_104_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13495_ (.CLK(clknet_leaf_105_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13496_ (.CLK(clknet_leaf_102_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13497_ (.CLK(clknet_leaf_103_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13498_ (.CLK(clknet_leaf_103_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13499_ (.CLK(clknet_leaf_103_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13500_ (.CLK(clknet_leaf_103_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13501_ (.CLK(clknet_leaf_123_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13502_ (.CLK(clknet_leaf_123_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13503_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13504_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13505_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13506_ (.CLK(clknet_leaf_123_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13507_ (.CLK(clknet_leaf_124_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13508_ (.CLK(clknet_leaf_123_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13509_ (.CLK(clknet_leaf_123_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13510_ (.CLK(clknet_leaf_105_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij._00_[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._23_[32] ));
 sky130_fd_sc_hd__dfxtp_1 _13511_ (.CLK(clknet_leaf_92_clk),
    .D(\sa_inst.sak._03_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._19_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13512_ (.CLK(clknet_leaf_84_clk),
    .D(\sa_inst.sak._03_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._19_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13513_ (.CLK(clknet_leaf_84_clk),
    .D(\sa_inst.sak._03_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._19_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13514_ (.CLK(clknet_leaf_84_clk),
    .D(\sa_inst.sak._03_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._19_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13515_ (.CLK(clknet_leaf_87_clk),
    .D(\sa_inst.sak._03_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._19_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13516_ (.CLK(clknet_leaf_87_clk),
    .D(\sa_inst.sak._03_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._19_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13517_ (.CLK(clknet_leaf_87_clk),
    .D(\sa_inst.sak._03_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._19_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13518_ (.CLK(clknet_leaf_87_clk),
    .D(\sa_inst.sak._03_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._19_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13519_ (.CLK(clknet_leaf_87_clk),
    .D(\sa_inst.sak._03_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._19_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13520_ (.CLK(clknet_leaf_87_clk),
    .D(\sa_inst.sak._03_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._19_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13521_ (.CLK(clknet_leaf_105_clk),
    .D(\sa_inst.sak._03_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._19_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13522_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak._04_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._20_ ));
 sky130_fd_sc_hd__dfrtp_1 _13523_ (.CLK(clknet_leaf_62_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[0] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13524_ (.CLK(clknet_leaf_60_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[1] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13525_ (.CLK(clknet_leaf_62_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[2] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13526_ (.CLK(clknet_leaf_64_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[3] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13527_ (.CLK(clknet_leaf_64_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[4] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13528_ (.CLK(clknet_leaf_64_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[5] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[5] ));
 sky130_fd_sc_hd__dfrtp_2 _13529_ (.CLK(clknet_leaf_65_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[6] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[6] ));
 sky130_fd_sc_hd__dfrtp_2 _13530_ (.CLK(clknet_leaf_65_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[7] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[7] ));
 sky130_fd_sc_hd__dfrtp_2 _13531_ (.CLK(clknet_leaf_67_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[8] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[8] ));
 sky130_fd_sc_hd__dfrtp_2 _13532_ (.CLK(clknet_leaf_67_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[9] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[9] ));
 sky130_fd_sc_hd__dfrtp_2 _13533_ (.CLK(clknet_leaf_65_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[10] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13534_ (.CLK(clknet_leaf_65_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[11] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13535_ (.CLK(clknet_leaf_68_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[12] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13536_ (.CLK(clknet_leaf_23_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[13] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[13] ));
 sky130_fd_sc_hd__dfrtp_2 _13537_ (.CLK(clknet_leaf_22_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[14] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[14] ));
 sky130_fd_sc_hd__dfrtp_2 _13538_ (.CLK(clknet_leaf_23_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[15] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[15] ));
 sky130_fd_sc_hd__dfrtp_2 _13539_ (.CLK(clknet_leaf_23_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[16] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[16] ));
 sky130_fd_sc_hd__dfrtp_2 _13540_ (.CLK(clknet_leaf_23_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[17] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13541_ (.CLK(clknet_leaf_23_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[18] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[18] ));
 sky130_fd_sc_hd__dfrtp_2 _13542_ (.CLK(clknet_leaf_23_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[19] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[19] ));
 sky130_fd_sc_hd__dfrtp_2 _13543_ (.CLK(clknet_leaf_24_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[20] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[20] ));
 sky130_fd_sc_hd__dfrtp_2 _13544_ (.CLK(clknet_leaf_21_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[21] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[21] ));
 sky130_fd_sc_hd__dfrtp_2 _13545_ (.CLK(clknet_leaf_19_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[22] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[22] ));
 sky130_fd_sc_hd__dfrtp_2 _13546_ (.CLK(clknet_leaf_19_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[23] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[23] ));
 sky130_fd_sc_hd__dfrtp_4 _13547_ (.CLK(clknet_leaf_20_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[24] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[24] ));
 sky130_fd_sc_hd__dfrtp_4 _13548_ (.CLK(clknet_leaf_20_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[25] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[25] ));
 sky130_fd_sc_hd__dfrtp_4 _13549_ (.CLK(clknet_leaf_164_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[26] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[26] ));
 sky130_fd_sc_hd__dfrtp_4 _13550_ (.CLK(clknet_leaf_163_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[27] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[27] ));
 sky130_fd_sc_hd__dfrtp_4 _13551_ (.CLK(clknet_leaf_21_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[28] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[28] ));
 sky130_fd_sc_hd__dfrtp_4 _13552_ (.CLK(clknet_leaf_21_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[29] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[29] ));
 sky130_fd_sc_hd__dfrtp_4 _13553_ (.CLK(clknet_leaf_22_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[30] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[30] ));
 sky130_fd_sc_hd__dfrtp_2 _13554_ (.CLK(clknet_leaf_22_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._24_[31] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._10_[31] ));
 sky130_fd_sc_hd__dfrtp_1 _13555_ (.CLK(clknet_leaf_69_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij.s3fdp_inst._20_ ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:1.pe_ij._02_ ));
 sky130_fd_sc_hd__dfxtp_1 _13556_ (.CLK(clknet_leaf_23_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13557_ (.CLK(clknet_leaf_23_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13558_ (.CLK(clknet_leaf_23_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13559_ (.CLK(clknet_leaf_26_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13560_ (.CLK(clknet_leaf_24_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13561_ (.CLK(clknet_leaf_26_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13562_ (.CLK(clknet_leaf_24_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13563_ (.CLK(clknet_leaf_19_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13564_ (.CLK(clknet_leaf_25_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13565_ (.CLK(clknet_leaf_26_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13566_ (.CLK(clknet_leaf_25_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13567_ (.CLK(clknet_leaf_25_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13568_ (.CLK(clknet_leaf_25_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13569_ (.CLK(clknet_leaf_18_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13570_ (.CLK(clknet_leaf_12_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13571_ (.CLK(clknet_leaf_13_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13572_ (.CLK(clknet_leaf_18_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13573_ (.CLK(clknet_leaf_18_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13574_ (.CLK(clknet_leaf_25_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13575_ (.CLK(clknet_leaf_13_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13576_ (.CLK(clknet_leaf_13_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13577_ (.CLK(clknet_leaf_13_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13578_ (.CLK(clknet_leaf_13_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13579_ (.CLK(clknet_leaf_13_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13580_ (.CLK(clknet_leaf_5_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13581_ (.CLK(clknet_leaf_5_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13582_ (.CLK(clknet_leaf_5_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13583_ (.CLK(clknet_leaf_14_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13584_ (.CLK(clknet_leaf_14_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13585_ (.CLK(clknet_leaf_14_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13586_ (.CLK(clknet_leaf_14_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[30] ));
 sky130_fd_sc_hd__dfxtp_2 _13587_ (.CLK(clknet_leaf_19_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13588_ (.CLK(clknet_leaf_163_clk),
    .D(\sa_inst.sak.rows:3.cols:1.pe_ij._00_[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[32] ));
 sky130_fd_sc_hd__dfrtp_1 _13589_ (.CLK(clknet_leaf_84_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[0] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13590_ (.CLK(clknet_leaf_75_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[1] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13591_ (.CLK(clknet_leaf_74_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[2] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13592_ (.CLK(clknet_leaf_74_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[3] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13593_ (.CLK(clknet_leaf_74_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[4] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13594_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[5] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[5] ));
 sky130_fd_sc_hd__dfrtp_4 _13595_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[6] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13596_ (.CLK(clknet_leaf_73_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[7] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13597_ (.CLK(clknet_leaf_106_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[8] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13598_ (.CLK(clknet_leaf_106_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[9] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13599_ (.CLK(clknet_leaf_107_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[10] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13600_ (.CLK(clknet_leaf_107_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[11] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13601_ (.CLK(clknet_leaf_107_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[12] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13602_ (.CLK(clknet_leaf_104_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[13] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13603_ (.CLK(clknet_leaf_108_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[14] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13604_ (.CLK(clknet_leaf_108_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[15] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[15] ));
 sky130_fd_sc_hd__dfrtp_2 _13605_ (.CLK(clknet_leaf_109_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[16] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[16] ));
 sky130_fd_sc_hd__dfrtp_2 _13606_ (.CLK(clknet_leaf_111_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[17] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[17] ));
 sky130_fd_sc_hd__dfrtp_2 _13607_ (.CLK(clknet_leaf_110_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[18] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[18] ));
 sky130_fd_sc_hd__dfrtp_2 _13608_ (.CLK(clknet_leaf_110_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[19] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[19] ));
 sky130_fd_sc_hd__dfrtp_2 _13609_ (.CLK(clknet_leaf_110_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[20] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[20] ));
 sky130_fd_sc_hd__dfrtp_2 _13610_ (.CLK(clknet_leaf_110_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[21] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[21] ));
 sky130_fd_sc_hd__dfrtp_2 _13611_ (.CLK(clknet_leaf_116_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[22] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[22] ));
 sky130_fd_sc_hd__dfrtp_2 _13612_ (.CLK(clknet_leaf_115_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[23] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[23] ));
 sky130_fd_sc_hd__dfrtp_2 _13613_ (.CLK(clknet_leaf_117_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[24] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[24] ));
 sky130_fd_sc_hd__dfrtp_2 _13614_ (.CLK(clknet_leaf_117_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[25] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13615_ (.CLK(clknet_leaf_115_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[26] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13616_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[27] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[27] ));
 sky130_fd_sc_hd__dfrtp_1 _13617_ (.CLK(clknet_leaf_114_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[28] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[28] ));
 sky130_fd_sc_hd__dfrtp_1 _13618_ (.CLK(clknet_leaf_115_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[29] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[29] ));
 sky130_fd_sc_hd__dfrtp_1 _13619_ (.CLK(clknet_leaf_115_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[30] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[30] ));
 sky130_fd_sc_hd__dfrtp_1 _13620_ (.CLK(clknet_leaf_116_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._24_[31] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._10_[31] ));
 sky130_fd_sc_hd__dfrtp_1 _13621_ (.CLK(clknet_leaf_107_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij.s3fdp_inst._20_ ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:2.pe_ij._02_ ));
 sky130_fd_sc_hd__dfxtp_1 _13622_ (.CLK(clknet_leaf_116_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[33] ));
 sky130_fd_sc_hd__dfxtp_1 _13623_ (.CLK(clknet_leaf_117_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[34] ));
 sky130_fd_sc_hd__dfxtp_1 _13624_ (.CLK(clknet_leaf_117_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[35] ));
 sky130_fd_sc_hd__dfxtp_1 _13625_ (.CLK(clknet_leaf_117_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[36] ));
 sky130_fd_sc_hd__dfxtp_1 _13626_ (.CLK(clknet_leaf_122_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[37] ));
 sky130_fd_sc_hd__dfxtp_1 _13627_ (.CLK(clknet_leaf_117_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[38] ));
 sky130_fd_sc_hd__dfxtp_1 _13628_ (.CLK(clknet_leaf_117_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[39] ));
 sky130_fd_sc_hd__dfxtp_1 _13629_ (.CLK(clknet_leaf_119_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[40] ));
 sky130_fd_sc_hd__dfxtp_1 _13630_ (.CLK(clknet_leaf_119_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[41] ));
 sky130_fd_sc_hd__dfxtp_1 _13631_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[42] ));
 sky130_fd_sc_hd__dfxtp_1 _13632_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[43] ));
 sky130_fd_sc_hd__dfxtp_1 _13633_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[44] ));
 sky130_fd_sc_hd__dfxtp_1 _13634_ (.CLK(clknet_leaf_120_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[45] ));
 sky130_fd_sc_hd__dfxtp_1 _13635_ (.CLK(clknet_leaf_117_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[46] ));
 sky130_fd_sc_hd__dfxtp_1 _13636_ (.CLK(clknet_leaf_118_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[47] ));
 sky130_fd_sc_hd__dfxtp_1 _13637_ (.CLK(clknet_leaf_118_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[48] ));
 sky130_fd_sc_hd__dfxtp_1 _13638_ (.CLK(clknet_leaf_118_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[49] ));
 sky130_fd_sc_hd__dfxtp_1 _13639_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[50] ));
 sky130_fd_sc_hd__dfxtp_1 _13640_ (.CLK(clknet_leaf_118_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[51] ));
 sky130_fd_sc_hd__dfxtp_1 _13641_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[52] ));
 sky130_fd_sc_hd__dfxtp_1 _13642_ (.CLK(clknet_leaf_118_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[53] ));
 sky130_fd_sc_hd__dfxtp_1 _13643_ (.CLK(clknet_leaf_118_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[54] ));
 sky130_fd_sc_hd__dfxtp_1 _13644_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[55] ));
 sky130_fd_sc_hd__dfxtp_1 _13645_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[56] ));
 sky130_fd_sc_hd__dfxtp_1 _13646_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[57] ));
 sky130_fd_sc_hd__dfxtp_1 _13647_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[58] ));
 sky130_fd_sc_hd__dfxtp_1 _13648_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[59] ));
 sky130_fd_sc_hd__dfxtp_1 _13649_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[60] ));
 sky130_fd_sc_hd__dfxtp_1 _13650_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[61] ));
 sky130_fd_sc_hd__dfxtp_1 _13651_ (.CLK(clknet_leaf_157_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[62] ));
 sky130_fd_sc_hd__dfxtp_1 _13652_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[63] ));
 sky130_fd_sc_hd__dfxtp_2 _13653_ (.CLK(clknet_leaf_118_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[64] ));
 sky130_fd_sc_hd__dfxtp_1 _13654_ (.CLK(clknet_leaf_143_clk),
    .D(\sa_inst.sak.rows:3.cols:2.pe_ij._00_[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[65] ));
 sky130_fd_sc_hd__dfxtp_1 _13655_ (.CLK(clknet_leaf_77_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13656_ (.CLK(clknet_leaf_77_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13657_ (.CLK(clknet_leaf_77_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13658_ (.CLK(clknet_leaf_78_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13659_ (.CLK(clknet_leaf_58_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13660_ (.CLK(clknet_leaf_58_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13661_ (.CLK(clknet_leaf_58_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13662_ (.CLK(clknet_leaf_58_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13663_ (.CLK(clknet_leaf_58_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13664_ (.CLK(clknet_leaf_58_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13665_ (.CLK(clknet_leaf_58_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13666_ (.CLK(clknet_leaf_58_clk),
    .D(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13667_ (.CLK(clknet_leaf_91_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[0] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13668_ (.CLK(clknet_leaf_91_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[1] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13669_ (.CLK(clknet_leaf_91_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[2] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13670_ (.CLK(clknet_leaf_90_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[3] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13671_ (.CLK(clknet_leaf_90_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[4] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13672_ (.CLK(clknet_leaf_90_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[5] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13673_ (.CLK(clknet_leaf_90_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[6] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13674_ (.CLK(clknet_leaf_97_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[7] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13675_ (.CLK(clknet_leaf_91_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[8] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13676_ (.CLK(clknet_leaf_95_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[9] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13677_ (.CLK(clknet_leaf_96_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[10] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13678_ (.CLK(clknet_leaf_97_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[11] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13679_ (.CLK(clknet_leaf_97_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[12] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13680_ (.CLK(clknet_leaf_97_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[13] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13681_ (.CLK(clknet_leaf_96_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[14] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13682_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[15] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13683_ (.CLK(clknet_leaf_102_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[16] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13684_ (.CLK(clknet_leaf_102_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[17] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13685_ (.CLK(clknet_leaf_105_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[18] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13686_ (.CLK(clknet_leaf_102_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[19] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13687_ (.CLK(clknet_leaf_103_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[20] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13688_ (.CLK(clknet_leaf_103_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[21] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13689_ (.CLK(clknet_leaf_103_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[22] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13690_ (.CLK(clknet_leaf_123_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[23] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[23] ));
 sky130_fd_sc_hd__dfrtp_2 _13691_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[24] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13692_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[25] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13693_ (.CLK(clknet_leaf_124_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[26] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13694_ (.CLK(clknet_leaf_124_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[27] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[27] ));
 sky130_fd_sc_hd__dfrtp_1 _13695_ (.CLK(clknet_leaf_121_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[28] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[28] ));
 sky130_fd_sc_hd__dfrtp_1 _13696_ (.CLK(clknet_leaf_124_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[29] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[29] ));
 sky130_fd_sc_hd__dfrtp_1 _13697_ (.CLK(clknet_leaf_124_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[30] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[30] ));
 sky130_fd_sc_hd__dfrtp_1 _13698_ (.CLK(clknet_leaf_123_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._24_[31] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._10_[31] ));
 sky130_fd_sc_hd__dfrtp_1 _13699_ (.CLK(clknet_leaf_94_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._20_ ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._02_ ));
 sky130_fd_sc_hd__dfxtp_2 _13700_ (.CLK(clknet_leaf_103_clk),
    .D(\sa_inst.EOB_Q_o ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij._01_ ));
 sky130_fd_sc_hd__dfxtp_1 _13701_ (.CLK(clknet_leaf_93_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._17_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._26_ ));
 sky130_fd_sc_hd__dfxtp_1 _13702_ (.CLK(clknet_leaf_93_clk),
    .D(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._25_ ));
 sky130_fd_sc_hd__dfxtp_1 _13703_ (.CLK(clknet_leaf_91_clk),
    .D(\sa_inst.sak._19_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._22_ ));
 sky130_fd_sc_hd__dfxtp_1 _13704_ (.CLK(clknet_leaf_105_clk),
    .D(\sa_inst.sak._19_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst._11_ ));
 sky130_fd_sc_hd__dfxtp_2 _13705_ (.CLK(clknet_leaf_57_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j._12_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._06_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13706_ (.CLK(clknet_leaf_56_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j._12_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._06_[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13707_ (.CLK(clknet_leaf_56_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j._12_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._06_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13708_ (.CLK(clknet_leaf_56_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j._12_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._06_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13709_ (.CLK(clknet_leaf_89_clk),
    .D(\sa_inst.sak._19_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13710_ (.CLK(clknet_leaf_92_clk),
    .D(\sa_inst.sak._19_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13711_ (.CLK(clknet_leaf_91_clk),
    .D(\sa_inst.sak._19_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._0_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13712_ (.CLK(clknet_leaf_86_clk),
    .D(_00135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13713_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[66] ));
 sky130_fd_sc_hd__dfxtp_1 _13714_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[67] ));
 sky130_fd_sc_hd__dfxtp_1 _13715_ (.CLK(clknet_leaf_99_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[68] ));
 sky130_fd_sc_hd__dfxtp_1 _13716_ (.CLK(clknet_leaf_99_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[69] ));
 sky130_fd_sc_hd__dfxtp_1 _13717_ (.CLK(clknet_leaf_99_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[70] ));
 sky130_fd_sc_hd__dfxtp_1 _13718_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[71] ));
 sky130_fd_sc_hd__dfxtp_1 _13719_ (.CLK(clknet_leaf_99_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[72] ));
 sky130_fd_sc_hd__dfxtp_1 _13720_ (.CLK(clknet_leaf_94_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[73] ));
 sky130_fd_sc_hd__dfxtp_1 _13721_ (.CLK(clknet_leaf_95_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[74] ));
 sky130_fd_sc_hd__dfxtp_1 _13722_ (.CLK(clknet_leaf_94_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[75] ));
 sky130_fd_sc_hd__dfxtp_1 _13723_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[76] ));
 sky130_fd_sc_hd__dfxtp_1 _13724_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[77] ));
 sky130_fd_sc_hd__dfxtp_1 _13725_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[78] ));
 sky130_fd_sc_hd__dfxtp_1 _13726_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[79] ));
 sky130_fd_sc_hd__dfxtp_1 _13727_ (.CLK(clknet_leaf_98_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[80] ));
 sky130_fd_sc_hd__dfxtp_1 _13728_ (.CLK(clknet_leaf_101_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[81] ));
 sky130_fd_sc_hd__dfxtp_1 _13729_ (.CLK(clknet_leaf_101_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[82] ));
 sky130_fd_sc_hd__dfxtp_1 _13730_ (.CLK(clknet_leaf_101_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[83] ));
 sky130_fd_sc_hd__dfxtp_1 _13731_ (.CLK(clknet_leaf_101_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[84] ));
 sky130_fd_sc_hd__dfxtp_1 _13732_ (.CLK(clknet_leaf_101_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[85] ));
 sky130_fd_sc_hd__dfxtp_1 _13733_ (.CLK(clknet_leaf_101_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[86] ));
 sky130_fd_sc_hd__dfxtp_1 _13734_ (.CLK(clknet_leaf_101_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[87] ));
 sky130_fd_sc_hd__dfxtp_1 _13735_ (.CLK(clknet_leaf_101_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[88] ));
 sky130_fd_sc_hd__dfxtp_1 _13736_ (.CLK(clknet_leaf_101_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[89] ));
 sky130_fd_sc_hd__dfxtp_1 _13737_ (.CLK(clknet_leaf_125_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[90] ));
 sky130_fd_sc_hd__dfxtp_1 _13738_ (.CLK(clknet_leaf_127_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[91] ));
 sky130_fd_sc_hd__dfxtp_1 _13739_ (.CLK(clknet_leaf_124_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[92] ));
 sky130_fd_sc_hd__dfxtp_1 _13740_ (.CLK(clknet_leaf_124_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[93] ));
 sky130_fd_sc_hd__dfxtp_1 _13741_ (.CLK(clknet_leaf_124_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[94] ));
 sky130_fd_sc_hd__dfxtp_1 _13742_ (.CLK(clknet_leaf_124_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[95] ));
 sky130_fd_sc_hd__dfxtp_1 _13743_ (.CLK(clknet_leaf_125_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[96] ));
 sky130_fd_sc_hd__dfxtp_1 _13744_ (.CLK(clknet_leaf_125_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[97] ));
 sky130_fd_sc_hd__dfxtp_1 _13745_ (.CLK(clknet_leaf_131_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij._00_[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._12_[98] ));
 sky130_fd_sc_hd__dfxtp_4 _13746_ (.CLK(clknet_leaf_83_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j._15_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._07_[0] ));
 sky130_fd_sc_hd__dfxtp_2 _13747_ (.CLK(clknet_leaf_83_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j._15_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:3.a2s3_j._23_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13748_ (.CLK(clknet_leaf_84_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j._15_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:3.a2s3_j._23_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13749_ (.CLK(clknet_leaf_83_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j._15_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:3.a2s3_j._23_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13750_ (.CLK(clknet_leaf_47_clk),
    .D(_00136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._05_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13751_ (.CLK(clknet_leaf_53_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j._07_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:2.a2s3_j._19_ ));
 sky130_fd_sc_hd__dfxtp_2 _13752_ (.CLK(clknet_leaf_53_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j._17_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._06_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13753_ (.CLK(clknet_leaf_53_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:2.a2s3_j._17_ ));
 sky130_fd_sc_hd__dfxtp_1 _13754_ (.CLK(clknet_leaf_55_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._01_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._10_ ));
 sky130_fd_sc_hd__dfxtp_1 _13755_ (.CLK(clknet_leaf_182_clk),
    .D(_00137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13756_ (.CLK(clknet_leaf_187_clk),
    .D(_00138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13757_ (.CLK(clknet_leaf_179_clk),
    .D(_00139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13758_ (.CLK(clknet_leaf_179_clk),
    .D(_00140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13759_ (.CLK(clknet_leaf_178_clk),
    .D(_00141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13760_ (.CLK(clknet_leaf_159_clk),
    .D(_00142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13761_ (.CLK(clknet_leaf_154_clk),
    .D(_00143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13762_ (.CLK(clknet_leaf_159_clk),
    .D(_00144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13763_ (.CLK(clknet_leaf_159_clk),
    .D(_00145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13764_ (.CLK(clknet_leaf_155_clk),
    .D(_00146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13765_ (.CLK(clknet_leaf_150_clk),
    .D(_00147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13766_ (.CLK(clknet_leaf_149_clk),
    .D(_00148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13767_ (.CLK(clknet_leaf_148_clk),
    .D(_00149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13768_ (.CLK(clknet_leaf_147_clk),
    .D(_00150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13769_ (.CLK(clknet_leaf_148_clk),
    .D(_00151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13770_ (.CLK(clknet_leaf_3_clk),
    .D(_00152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13771_ (.CLK(clknet_leaf_4_clk),
    .D(_00153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13772_ (.CLK(clknet_leaf_5_clk),
    .D(_00154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13773_ (.CLK(clknet_leaf_6_clk),
    .D(_00155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13774_ (.CLK(clknet_leaf_1_clk),
    .D(_00156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13775_ (.CLK(clknet_leaf_190_clk),
    .D(_00157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13776_ (.CLK(clknet_leaf_190_clk),
    .D(_00158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13777_ (.CLK(clknet_leaf_188_clk),
    .D(_00159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13778_ (.CLK(clknet_leaf_189_clk),
    .D(_00160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13779_ (.CLK(clknet_leaf_53_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j._15_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._05_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13780_ (.CLK(clknet_leaf_52_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j._15_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:1.a2s3_j._23_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13781_ (.CLK(clknet_leaf_52_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j._15_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:1.a2s3_j._23_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13782_ (.CLK(clknet_leaf_52_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j._15_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:1.a2s3_j._23_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13783_ (.CLK(clknet_leaf_99_clk),
    .D(_00161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13784_ (.CLK(clknet_leaf_100_clk),
    .D(_00162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13785_ (.CLK(clknet_leaf_100_clk),
    .D(_00163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13786_ (.CLK(clknet_leaf_99_clk),
    .D(_00164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13787_ (.CLK(clknet_leaf_99_clk),
    .D(_00165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13788_ (.CLK(clknet_leaf_99_clk),
    .D(_00166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13789_ (.CLK(clknet_leaf_99_clk),
    .D(_00167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13790_ (.CLK(clknet_leaf_99_clk),
    .D(_00168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13791_ (.CLK(clknet_leaf_125_clk),
    .D(_00169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13792_ (.CLK(clknet_leaf_99_clk),
    .D(_00170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13793_ (.CLK(clknet_leaf_99_clk),
    .D(_00171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13794_ (.CLK(clknet_leaf_100_clk),
    .D(_00172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13795_ (.CLK(clknet_leaf_125_clk),
    .D(_00173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13796_ (.CLK(clknet_leaf_100_clk),
    .D(_00174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13797_ (.CLK(clknet_leaf_100_clk),
    .D(_00175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13798_ (.CLK(clknet_leaf_100_clk),
    .D(_00176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13799_ (.CLK(clknet_leaf_99_clk),
    .D(_00177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13800_ (.CLK(clknet_leaf_100_clk),
    .D(_00178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13801_ (.CLK(clknet_leaf_100_clk),
    .D(_00179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13802_ (.CLK(clknet_leaf_100_clk),
    .D(_00180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13803_ (.CLK(clknet_leaf_125_clk),
    .D(_00181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13804_ (.CLK(clknet_leaf_125_clk),
    .D(_00182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13805_ (.CLK(clknet_leaf_101_clk),
    .D(_00183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13806_ (.CLK(clknet_leaf_125_clk),
    .D(_00184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13807_ (.CLK(clknet_leaf_124_clk),
    .D(_00185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13808_ (.CLK(clknet_leaf_124_clk),
    .D(_00186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13809_ (.CLK(clknet_leaf_124_clk),
    .D(_00187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13810_ (.CLK(clknet_leaf_124_clk),
    .D(_00188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13811_ (.CLK(clknet_leaf_124_clk),
    .D(_00189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13812_ (.CLK(clknet_leaf_125_clk),
    .D(_00190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13813_ (.CLK(clknet_leaf_125_clk),
    .D(_00191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._66_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13814_ (.CLK(clknet_leaf_52_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j._14_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:1.a2s3_j._15_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13815_ (.CLK(clknet_leaf_53_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j._19_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._05_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13816_ (.CLK(clknet_leaf_53_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j._07_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:1.a2s3_j._19_ ));
 sky130_fd_sc_hd__dfxtp_1 _13817_ (.CLK(clknet_leaf_61_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j._17_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._05_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13818_ (.CLK(clknet_leaf_61_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:1.a2s3_j._17_ ));
 sky130_fd_sc_hd__dfxtp_1 _13819_ (.CLK(clknet_leaf_181_clk),
    .D(_00192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13820_ (.CLK(clknet_leaf_188_clk),
    .D(_00193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13821_ (.CLK(clknet_leaf_181_clk),
    .D(_00194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13822_ (.CLK(clknet_leaf_181_clk),
    .D(_00195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13823_ (.CLK(clknet_leaf_181_clk),
    .D(_00196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13824_ (.CLK(clknet_leaf_167_clk),
    .D(_00197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13825_ (.CLK(clknet_leaf_173_clk),
    .D(_00198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13826_ (.CLK(clknet_leaf_160_clk),
    .D(_00199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13827_ (.CLK(clknet_leaf_174_clk),
    .D(_00200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13828_ (.CLK(clknet_leaf_154_clk),
    .D(_00201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13829_ (.CLK(clknet_leaf_150_clk),
    .D(_00202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13830_ (.CLK(clknet_leaf_150_clk),
    .D(_00203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13831_ (.CLK(clknet_leaf_150_clk),
    .D(_00204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13832_ (.CLK(clknet_leaf_178_clk),
    .D(_00205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13833_ (.CLK(clknet_leaf_178_clk),
    .D(_00206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13834_ (.CLK(clknet_leaf_5_clk),
    .D(_00207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13835_ (.CLK(clknet_leaf_4_clk),
    .D(_00208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13836_ (.CLK(clknet_leaf_6_clk),
    .D(_00209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13837_ (.CLK(clknet_leaf_6_clk),
    .D(_00210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13838_ (.CLK(clknet_leaf_1_clk),
    .D(_00211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13839_ (.CLK(clknet_leaf_190_clk),
    .D(_00212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13840_ (.CLK(clknet_leaf_190_clk),
    .D(_00213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13841_ (.CLK(clknet_leaf_188_clk),
    .D(_00214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13842_ (.CLK(clknet_leaf_190_clk),
    .D(_00215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[14][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13843_ (.CLK(clknet_leaf_125_clk),
    .D(\sa_inst._12_[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._00_ ));
 sky130_fd_sc_hd__dfxtp_1 _13844_ (.CLK(clknet_leaf_130_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._27_ ));
 sky130_fd_sc_hd__dfxtp_1 _13845_ (.CLK(clknet_leaf_132_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._25_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._26_ ));
 sky130_fd_sc_hd__dfxtp_1 _13846_ (.CLK(clknet_leaf_130_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._24_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._25_ ));
 sky130_fd_sc_hd__dfxtp_1 _13847_ (.CLK(clknet_leaf_120_clk),
    .D(_00216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13848_ (.CLK(clknet_leaf_120_clk),
    .D(_00217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13849_ (.CLK(clknet_leaf_120_clk),
    .D(_00218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13850_ (.CLK(clknet_leaf_120_clk),
    .D(_00219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13851_ (.CLK(clknet_leaf_120_clk),
    .D(_00220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13852_ (.CLK(clknet_leaf_120_clk),
    .D(_00221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13853_ (.CLK(clknet_leaf_120_clk),
    .D(_00222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13854_ (.CLK(clknet_leaf_120_clk),
    .D(_00223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13855_ (.CLK(clknet_leaf_121_clk),
    .D(_00224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13856_ (.CLK(clknet_leaf_120_clk),
    .D(_00225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13857_ (.CLK(clknet_leaf_131_clk),
    .D(_00226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13858_ (.CLK(clknet_leaf_120_clk),
    .D(_00227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13859_ (.CLK(clknet_leaf_157_clk),
    .D(_00228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13860_ (.CLK(clknet_leaf_157_clk),
    .D(_00229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13861_ (.CLK(clknet_leaf_156_clk),
    .D(_00230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13862_ (.CLK(clknet_leaf_119_clk),
    .D(_00231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13863_ (.CLK(clknet_leaf_119_clk),
    .D(_00232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13864_ (.CLK(clknet_leaf_119_clk),
    .D(_00233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13865_ (.CLK(clknet_leaf_119_clk),
    .D(_00234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13866_ (.CLK(clknet_leaf_119_clk),
    .D(_00235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13867_ (.CLK(clknet_leaf_119_clk),
    .D(_00236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13868_ (.CLK(clknet_leaf_119_clk),
    .D(_00237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13869_ (.CLK(clknet_leaf_119_clk),
    .D(_00238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13870_ (.CLK(clknet_leaf_157_clk),
    .D(_00239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13871_ (.CLK(clknet_leaf_157_clk),
    .D(_00240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13872_ (.CLK(clknet_leaf_157_clk),
    .D(_00241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13873_ (.CLK(clknet_leaf_157_clk),
    .D(_00242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13874_ (.CLK(clknet_leaf_157_clk),
    .D(_00243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13875_ (.CLK(clknet_leaf_157_clk),
    .D(_00244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13876_ (.CLK(clknet_leaf_157_clk),
    .D(_00245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13877_ (.CLK(clknet_leaf_157_clk),
    .D(_00246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._66_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13878_ (.CLK(clknet_leaf_156_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._21_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._23_ ));
 sky130_fd_sc_hd__dfxtp_1 _13879_ (.CLK(clknet_leaf_156_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._20_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._21_ ));
 sky130_fd_sc_hd__dfxtp_1 _13880_ (.CLK(clknet_leaf_156_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._19_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._20_ ));
 sky130_fd_sc_hd__dfxtp_1 _13881_ (.CLK(clknet_leaf_156_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._18_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._19_ ));
 sky130_fd_sc_hd__dfxtp_1 _13882_ (.CLK(clknet_leaf_156_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._17_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._18_ ));
 sky130_fd_sc_hd__dfxtp_1 _13883_ (.CLK(clknet_leaf_156_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._16_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._17_ ));
 sky130_fd_sc_hd__dfxtp_1 _13884_ (.CLK(clknet_leaf_157_clk),
    .D(\sa_inst._12_[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._16_ ));
 sky130_fd_sc_hd__dfxtp_2 _13885_ (.CLK(clknet_leaf_134_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._46_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._15_ ));
 sky130_fd_sc_hd__dfxtp_1 _13886_ (.CLK(clknet_leaf_134_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._13_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._14_ ));
 sky130_fd_sc_hd__dfxtp_1 _13887_ (.CLK(clknet_leaf_134_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._40_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._13_ ));
 sky130_fd_sc_hd__dfxtp_2 _13888_ (.CLK(clknet_leaf_135_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._08_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._09_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13889_ (.CLK(clknet_leaf_143_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._08_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._09_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13890_ (.CLK(clknet_leaf_156_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._08_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._09_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13891_ (.CLK(clknet_leaf_143_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._08_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._09_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13892_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._08_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._09_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13893_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._08_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._09_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13894_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._08_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._09_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13895_ (.CLK(clknet_leaf_135_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._07_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._08_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13896_ (.CLK(clknet_leaf_135_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._07_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._08_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13897_ (.CLK(clknet_leaf_156_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._07_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._08_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13898_ (.CLK(clknet_leaf_143_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._07_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._08_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13899_ (.CLK(clknet_leaf_143_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._07_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._08_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13900_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._07_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._08_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13901_ (.CLK(clknet_leaf_134_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._07_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._08_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13902_ (.CLK(clknet_leaf_135_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._40_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._07_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13903_ (.CLK(clknet_leaf_134_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._40_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._07_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13904_ (.CLK(clknet_leaf_143_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._40_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._07_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13905_ (.CLK(clknet_leaf_143_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._40_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._07_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13906_ (.CLK(clknet_leaf_143_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._40_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._07_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13907_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._40_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._07_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13908_ (.CLK(clknet_leaf_134_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._37_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._07_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13909_ (.CLK(clknet_leaf_131_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._31_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._06_ ));
 sky130_fd_sc_hd__dfxtp_1 _13910_ (.CLK(clknet_leaf_129_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._31_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._05_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13911_ (.CLK(clknet_leaf_129_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._31_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._05_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13912_ (.CLK(clknet_leaf_131_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._31_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._05_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13913_ (.CLK(clknet_leaf_131_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._31_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._05_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13914_ (.CLK(clknet_leaf_136_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._03_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._04_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13915_ (.CLK(clknet_leaf_136_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._02_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._03_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13916_ (.CLK(clknet_leaf_129_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._29_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._02_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13917_ (.CLK(clknet_leaf_130_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._29_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._02_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13918_ (.CLK(clknet_leaf_130_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._29_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._02_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13919_ (.CLK(clknet_leaf_130_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._29_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._02_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13920_ (.CLK(clknet_leaf_130_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._29_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._02_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13921_ (.CLK(clknet_leaf_130_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._29_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._02_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13922_ (.CLK(clknet_leaf_136_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._57_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._01_ ));
 sky130_fd_sc_hd__dfxtp_1 _13923_ (.CLK(clknet_leaf_135_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._56_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._57_ ));
 sky130_fd_sc_hd__dfxtp_1 _13924_ (.CLK(clknet_leaf_136_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._30_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._56_ ));
 sky130_fd_sc_hd__dfxtp_1 _13925_ (.CLK(clknet_leaf_135_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._54_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._55_ ));
 sky130_fd_sc_hd__dfxtp_1 _13926_ (.CLK(clknet_leaf_132_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._44_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._54_ ));
 sky130_fd_sc_hd__dfxtp_1 _13927_ (.CLK(clknet_leaf_130_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._33_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._44_ ));
 sky130_fd_sc_hd__dfxtp_1 _13928_ (.CLK(clknet_leaf_130_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._22_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._33_ ));
 sky130_fd_sc_hd__dfxtp_1 _13929_ (.CLK(clknet_leaf_131_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._11_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._22_ ));
 sky130_fd_sc_hd__dfxtp_1 _13930_ (.CLK(clknet_leaf_128_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._00_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._11_ ));
 sky130_fd_sc_hd__dfxtp_1 _13931_ (.CLK(clknet_leaf_131_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._23_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._33_ ));
 sky130_fd_sc_hd__dfxtp_1 _13932_ (.CLK(clknet_leaf_131_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._33_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._44_ ));
 sky130_fd_sc_hd__dfxtp_1 _13933_ (.CLK(clknet_leaf_131_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._44_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._55_ ));
 sky130_fd_sc_hd__dfxtp_1 _13934_ (.CLK(clknet_leaf_126_clk),
    .D(_00247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._05_ ));
 sky130_fd_sc_hd__dfxtp_1 _13935_ (.CLK(clknet_leaf_128_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._31_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._88_ ));
 sky130_fd_sc_hd__dfxtp_1 _13936_ (.CLK(clknet_leaf_131_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._88_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._01_ ));
 sky130_fd_sc_hd__dfxtp_1 _13937_ (.CLK(clknet_leaf_126_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13938_ (.CLK(clknet_leaf_128_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13939_ (.CLK(clknet_leaf_129_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13940_ (.CLK(clknet_leaf_127_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13941_ (.CLK(clknet_leaf_126_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13942_ (.CLK(clknet_leaf_128_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13943_ (.CLK(clknet_leaf_127_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13944_ (.CLK(clknet_leaf_126_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13945_ (.CLK(clknet_leaf_100_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13946_ (.CLK(clknet_leaf_126_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13947_ (.CLK(clknet_leaf_126_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13948_ (.CLK(clknet_leaf_126_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13949_ (.CLK(clknet_leaf_126_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13950_ (.CLK(clknet_leaf_126_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13951_ (.CLK(clknet_leaf_127_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13952_ (.CLK(clknet_leaf_127_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13953_ (.CLK(clknet_leaf_127_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13954_ (.CLK(clknet_leaf_128_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13955_ (.CLK(clknet_leaf_128_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13956_ (.CLK(clknet_leaf_127_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13957_ (.CLK(clknet_leaf_127_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13958_ (.CLK(clknet_leaf_127_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13959_ (.CLK(clknet_leaf_127_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._35_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._02_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13960_ (.CLK(clknet_leaf_132_clk),
    .D(_00248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._24_ ));
 sky130_fd_sc_hd__dfxtp_2 _13961_ (.CLK(clknet_leaf_127_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._42_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._06_ ));
 sky130_fd_sc_hd__dfxtp_1 _13962_ (.CLK(clknet_leaf_128_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._07_ ));
 sky130_fd_sc_hd__dfxtp_1 _13963_ (.CLK(clknet_leaf_127_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._48_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._08_ ));
 sky130_fd_sc_hd__dfxtp_1 _13964_ (.CLK(clknet_leaf_126_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._50_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._09_ ));
 sky130_fd_sc_hd__dfxtp_1 _13965_ (.CLK(clknet_leaf_131_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._56_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i._31_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13966_ (.CLK(clknet_leaf_129_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13967_ (.CLK(clknet_leaf_129_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13968_ (.CLK(clknet_leaf_129_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13969_ (.CLK(clknet_leaf_129_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13970_ (.CLK(clknet_leaf_128_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13971_ (.CLK(clknet_leaf_129_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13972_ (.CLK(clknet_leaf_128_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13973_ (.CLK(clknet_leaf_131_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13974_ (.CLK(clknet_leaf_131_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13975_ (.CLK(clknet_leaf_131_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._59_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._12_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13976_ (.CLK(clknet_leaf_129_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._67_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._13_ ));
 sky130_fd_sc_hd__dfxtp_1 _13977_ (.CLK(clknet_leaf_131_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._69_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._14_ ));
 sky130_fd_sc_hd__dfxtp_1 _13978_ (.CLK(clknet_leaf_129_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._74_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.lzoc_inst._15_ ));
 sky130_fd_sc_hd__dfxtp_1 _13979_ (.CLK(clknet_leaf_181_clk),
    .D(_00249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13980_ (.CLK(clknet_leaf_182_clk),
    .D(_00250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13981_ (.CLK(clknet_leaf_181_clk),
    .D(_00251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13982_ (.CLK(clknet_leaf_181_clk),
    .D(_00252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13983_ (.CLK(clknet_leaf_179_clk),
    .D(_00253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13984_ (.CLK(clknet_leaf_167_clk),
    .D(_00254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13985_ (.CLK(clknet_leaf_174_clk),
    .D(_00255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13986_ (.CLK(clknet_leaf_159_clk),
    .D(_00256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13987_ (.CLK(clknet_leaf_166_clk),
    .D(_00257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13988_ (.CLK(clknet_leaf_154_clk),
    .D(_00258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13989_ (.CLK(clknet_leaf_150_clk),
    .D(_00259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13990_ (.CLK(clknet_leaf_150_clk),
    .D(_00260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13991_ (.CLK(clknet_leaf_150_clk),
    .D(_00261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13992_ (.CLK(clknet_leaf_178_clk),
    .D(_00262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13993_ (.CLK(clknet_leaf_178_clk),
    .D(_00263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13994_ (.CLK(clknet_leaf_4_clk),
    .D(_00264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13995_ (.CLK(clknet_leaf_4_clk),
    .D(_00265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13996_ (.CLK(clknet_leaf_6_clk),
    .D(_00266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13997_ (.CLK(clknet_leaf_6_clk),
    .D(_00267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13998_ (.CLK(clknet_leaf_1_clk),
    .D(_00268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13999_ (.CLK(clknet_leaf_190_clk),
    .D(_00269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14000_ (.CLK(clknet_leaf_190_clk),
    .D(_00270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14001_ (.CLK(clknet_leaf_188_clk),
    .D(_00271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14002_ (.CLK(clknet_leaf_188_clk),
    .D(_00272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[13][23] ));
 sky130_fd_sc_hd__dfxtp_2 _14003_ (.CLK(clknet_leaf_78_clk),
    .D(\sa_inst.sak._07_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._13_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14004_ (.CLK(clknet_leaf_78_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w2_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14005_ (.CLK(clknet_leaf_78_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w3_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14006_ (.CLK(clknet_leaf_78_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w4_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14007_ (.CLK(clknet_leaf_78_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w5_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14008_ (.CLK(clknet_leaf_75_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w6_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14009_ (.CLK(clknet_leaf_75_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w7_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14010_ (.CLK(clknet_leaf_84_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w8_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14011_ (.CLK(clknet_leaf_75_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w9_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14012_ (.CLK(clknet_leaf_75_clk),
    .D(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_inst.bh33_w10_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:2.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14013_ (.CLK(clknet_leaf_181_clk),
    .D(_00273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14014_ (.CLK(clknet_leaf_181_clk),
    .D(_00274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14015_ (.CLK(clknet_leaf_181_clk),
    .D(_00275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14016_ (.CLK(clknet_leaf_178_clk),
    .D(_00276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14017_ (.CLK(clknet_leaf_178_clk),
    .D(_00277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14018_ (.CLK(clknet_leaf_166_clk),
    .D(_00278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14019_ (.CLK(clknet_leaf_174_clk),
    .D(_00279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14020_ (.CLK(clknet_leaf_159_clk),
    .D(_00280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14021_ (.CLK(clknet_leaf_160_clk),
    .D(_00281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14022_ (.CLK(clknet_leaf_154_clk),
    .D(_00282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14023_ (.CLK(clknet_leaf_150_clk),
    .D(_00283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14024_ (.CLK(clknet_leaf_150_clk),
    .D(_00284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14025_ (.CLK(clknet_leaf_150_clk),
    .D(_00285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14026_ (.CLK(clknet_leaf_150_clk),
    .D(_00286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14027_ (.CLK(clknet_leaf_151_clk),
    .D(_00287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14028_ (.CLK(clknet_leaf_4_clk),
    .D(_00288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14029_ (.CLK(clknet_leaf_15_clk),
    .D(_00289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14030_ (.CLK(clknet_leaf_5_clk),
    .D(_00290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14031_ (.CLK(clknet_leaf_6_clk),
    .D(_00291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14032_ (.CLK(clknet_leaf_1_clk),
    .D(_00292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14033_ (.CLK(clknet_leaf_190_clk),
    .D(_00293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14034_ (.CLK(clknet_leaf_190_clk),
    .D(_00294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14035_ (.CLK(clknet_leaf_188_clk),
    .D(_00295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14036_ (.CLK(clknet_leaf_188_clk),
    .D(_00296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14037_ (.CLK(clknet_leaf_135_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.rshift._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.rshift._11_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14038_ (.CLK(clknet_leaf_135_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._35_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.rshift._22_ ));
 sky130_fd_sc_hd__dfxtp_1 _14039_ (.CLK(clknet_leaf_136_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.rshift._04_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.rshift._25_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14040_ (.CLK(clknet_leaf_130_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.rshift._04_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.rshift._25_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14041_ (.CLK(clknet_leaf_135_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.rshift._04_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.rshift._25_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14042_ (.CLK(clknet_leaf_130_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.rshift._04_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.rshift._25_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14043_ (.CLK(clknet_leaf_135_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.rshift._10_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.rshift._26_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14044_ (.CLK(clknet_leaf_135_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.rshift._10_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.rshift._26_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14045_ (.CLK(clknet_leaf_135_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.rshift._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.rshift._27_ ));
 sky130_fd_sc_hd__dfxtp_1 _14046_ (.CLK(clknet_leaf_134_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.rshift._17_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.rshift._28_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14047_ (.CLK(clknet_leaf_136_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i.rshift._28_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.rshift._18_ ));
 sky130_fd_sc_hd__dfxtp_1 _14048_ (.CLK(clknet_leaf_134_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._35_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.rshift._00_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14049_ (.CLK(clknet_leaf_135_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._35_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.rshift._00_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14050_ (.CLK(clknet_leaf_135_clk),
    .D(\sa_inst.cols_l2a:3.l2a_i._35_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:3.l2a_i.rshift._00_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14051_ (.CLK(clknet_leaf_182_clk),
    .D(_00297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14052_ (.CLK(clknet_leaf_187_clk),
    .D(_00298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14053_ (.CLK(clknet_leaf_183_clk),
    .D(_00299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14054_ (.CLK(clknet_leaf_179_clk),
    .D(_00300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14055_ (.CLK(clknet_leaf_179_clk),
    .D(_00301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14056_ (.CLK(clknet_leaf_174_clk),
    .D(_00302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14057_ (.CLK(clknet_leaf_175_clk),
    .D(_00303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14058_ (.CLK(clknet_leaf_153_clk),
    .D(_00304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14059_ (.CLK(clknet_leaf_174_clk),
    .D(_00305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14060_ (.CLK(clknet_leaf_153_clk),
    .D(_00306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14061_ (.CLK(clknet_leaf_151_clk),
    .D(_00307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14062_ (.CLK(clknet_leaf_151_clk),
    .D(_00308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14063_ (.CLK(clknet_leaf_151_clk),
    .D(_00309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14064_ (.CLK(clknet_leaf_177_clk),
    .D(_00310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14065_ (.CLK(clknet_leaf_177_clk),
    .D(_00311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14066_ (.CLK(clknet_leaf_2_clk),
    .D(_00312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14067_ (.CLK(clknet_leaf_3_clk),
    .D(_00313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14068_ (.CLK(clknet_leaf_0_clk),
    .D(_00314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14069_ (.CLK(clknet_leaf_0_clk),
    .D(_00315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14070_ (.CLK(clknet_leaf_0_clk),
    .D(_00316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14071_ (.CLK(clknet_leaf_191_clk),
    .D(_00317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14072_ (.CLK(clknet_leaf_191_clk),
    .D(_00318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14073_ (.CLK(clknet_leaf_189_clk),
    .D(_00319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14074_ (.CLK(clknet_leaf_189_clk),
    .D(_00320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14075_ (.CLK(clknet_leaf_119_clk),
    .D(\sa_inst._12_[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._00_ ));
 sky130_fd_sc_hd__dfxtp_1 _14076_ (.CLK(clknet_leaf_145_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._27_ ));
 sky130_fd_sc_hd__dfxtp_1 _14077_ (.CLK(clknet_leaf_145_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._25_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._26_ ));
 sky130_fd_sc_hd__dfxtp_1 _14078_ (.CLK(clknet_leaf_145_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._24_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._25_ ));
 sky130_fd_sc_hd__dfxtp_1 _14079_ (.CLK(clknet_leaf_17_clk),
    .D(_00321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14080_ (.CLK(clknet_leaf_20_clk),
    .D(_00322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14081_ (.CLK(clknet_leaf_17_clk),
    .D(_00323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14082_ (.CLK(clknet_leaf_20_clk),
    .D(_00324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14083_ (.CLK(clknet_leaf_17_clk),
    .D(_00325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14084_ (.CLK(clknet_leaf_17_clk),
    .D(_00326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14085_ (.CLK(clknet_leaf_17_clk),
    .D(_00327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14086_ (.CLK(clknet_leaf_17_clk),
    .D(_00328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14087_ (.CLK(clknet_leaf_18_clk),
    .D(_00329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14088_ (.CLK(clknet_leaf_18_clk),
    .D(_00330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14089_ (.CLK(clknet_leaf_18_clk),
    .D(_00331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14090_ (.CLK(clknet_leaf_18_clk),
    .D(_00332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14091_ (.CLK(clknet_leaf_18_clk),
    .D(_00333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14092_ (.CLK(clknet_leaf_13_clk),
    .D(_00334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14093_ (.CLK(clknet_leaf_13_clk),
    .D(_00335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14094_ (.CLK(clknet_leaf_18_clk),
    .D(_00336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14095_ (.CLK(clknet_leaf_17_clk),
    .D(_00337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14096_ (.CLK(clknet_leaf_17_clk),
    .D(_00338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14097_ (.CLK(clknet_leaf_13_clk),
    .D(_00339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14098_ (.CLK(clknet_leaf_18_clk),
    .D(_00340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14099_ (.CLK(clknet_leaf_13_clk),
    .D(_00341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14100_ (.CLK(clknet_leaf_13_clk),
    .D(_00342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14101_ (.CLK(clknet_leaf_13_clk),
    .D(_00343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14102_ (.CLK(clknet_leaf_14_clk),
    .D(_00344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14103_ (.CLK(clknet_leaf_15_clk),
    .D(_00345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14104_ (.CLK(clknet_leaf_15_clk),
    .D(_00346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14105_ (.CLK(clknet_leaf_14_clk),
    .D(_00347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14106_ (.CLK(clknet_leaf_14_clk),
    .D(_00348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14107_ (.CLK(clknet_leaf_14_clk),
    .D(_00349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14108_ (.CLK(clknet_leaf_14_clk),
    .D(_00350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14109_ (.CLK(clknet_leaf_13_clk),
    .D(_00351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._66_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14110_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._21_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._23_ ));
 sky130_fd_sc_hd__dfxtp_1 _14111_ (.CLK(clknet_leaf_143_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._20_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._21_ ));
 sky130_fd_sc_hd__dfxtp_1 _14112_ (.CLK(clknet_leaf_143_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._19_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._20_ ));
 sky130_fd_sc_hd__dfxtp_1 _14113_ (.CLK(clknet_leaf_144_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._18_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._19_ ));
 sky130_fd_sc_hd__dfxtp_1 _14114_ (.CLK(clknet_leaf_143_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._17_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._18_ ));
 sky130_fd_sc_hd__dfxtp_1 _14115_ (.CLK(clknet_leaf_144_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._16_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._17_ ));
 sky130_fd_sc_hd__dfxtp_1 _14116_ (.CLK(clknet_leaf_144_clk),
    .D(\sa_inst._12_[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._16_ ));
 sky130_fd_sc_hd__dfxtp_1 _14117_ (.CLK(clknet_leaf_138_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._46_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._15_ ));
 sky130_fd_sc_hd__dfxtp_1 _14118_ (.CLK(clknet_leaf_138_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._13_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._14_ ));
 sky130_fd_sc_hd__dfxtp_1 _14119_ (.CLK(clknet_leaf_138_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._40_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._13_ ));
 sky130_fd_sc_hd__dfxtp_1 _14120_ (.CLK(clknet_leaf_139_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._08_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._09_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14121_ (.CLK(clknet_leaf_139_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._08_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._09_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14122_ (.CLK(clknet_leaf_138_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._08_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._09_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14123_ (.CLK(clknet_leaf_139_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._08_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._09_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14124_ (.CLK(clknet_leaf_147_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._08_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._09_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14125_ (.CLK(clknet_leaf_146_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._08_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._09_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14126_ (.CLK(clknet_leaf_138_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._08_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._09_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14127_ (.CLK(clknet_leaf_140_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._07_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._08_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14128_ (.CLK(clknet_leaf_139_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._07_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._08_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14129_ (.CLK(clknet_leaf_138_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._07_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._08_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14130_ (.CLK(clknet_leaf_139_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._07_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._08_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14131_ (.CLK(clknet_leaf_147_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._07_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._08_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14132_ (.CLK(clknet_leaf_147_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._07_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._08_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14133_ (.CLK(clknet_leaf_138_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._07_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._08_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14134_ (.CLK(clknet_leaf_139_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._40_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._07_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14135_ (.CLK(clknet_leaf_139_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._40_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._07_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14136_ (.CLK(clknet_leaf_138_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._40_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._07_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14137_ (.CLK(clknet_leaf_139_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._40_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._07_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14138_ (.CLK(clknet_leaf_147_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._40_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._07_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14139_ (.CLK(clknet_leaf_147_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._40_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._07_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14140_ (.CLK(clknet_leaf_138_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._37_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._07_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14141_ (.CLK(clknet_leaf_139_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._31_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._06_ ));
 sky130_fd_sc_hd__dfxtp_1 _14142_ (.CLK(clknet_leaf_137_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._31_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._05_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14143_ (.CLK(clknet_leaf_137_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._31_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._05_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14144_ (.CLK(clknet_leaf_139_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._31_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._05_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14145_ (.CLK(clknet_leaf_139_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._31_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._05_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14146_ (.CLK(clknet_leaf_137_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._03_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._04_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14147_ (.CLK(clknet_leaf_137_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._02_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._03_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14148_ (.CLK(clknet_leaf_140_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._29_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._02_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14149_ (.CLK(clknet_leaf_140_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._29_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._02_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14150_ (.CLK(clknet_leaf_140_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._29_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._02_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14151_ (.CLK(clknet_leaf_140_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._29_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._02_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14152_ (.CLK(clknet_leaf_140_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._29_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._02_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14153_ (.CLK(clknet_leaf_140_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._29_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._02_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14154_ (.CLK(clknet_leaf_137_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._57_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._01_ ));
 sky130_fd_sc_hd__dfxtp_1 _14155_ (.CLK(clknet_leaf_137_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._56_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._57_ ));
 sky130_fd_sc_hd__dfxtp_1 _14156_ (.CLK(clknet_leaf_141_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._30_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._56_ ));
 sky130_fd_sc_hd__dfxtp_1 _14157_ (.CLK(clknet_leaf_139_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._54_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._55_ ));
 sky130_fd_sc_hd__dfxtp_1 _14158_ (.CLK(clknet_leaf_139_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._44_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._54_ ));
 sky130_fd_sc_hd__dfxtp_1 _14159_ (.CLK(clknet_leaf_139_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._33_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._44_ ));
 sky130_fd_sc_hd__dfxtp_1 _14160_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._22_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._33_ ));
 sky130_fd_sc_hd__dfxtp_1 _14161_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._11_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._22_ ));
 sky130_fd_sc_hd__dfxtp_1 _14162_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._00_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._11_ ));
 sky130_fd_sc_hd__dfxtp_1 _14163_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._23_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._33_ ));
 sky130_fd_sc_hd__dfxtp_1 _14164_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._33_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._44_ ));
 sky130_fd_sc_hd__dfxtp_1 _14165_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._44_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._55_ ));
 sky130_fd_sc_hd__dfxtp_1 _14166_ (.CLK(clknet_leaf_132_clk),
    .D(_00352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._05_ ));
 sky130_fd_sc_hd__dfxtp_1 _14167_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._31_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._88_ ));
 sky130_fd_sc_hd__dfxtp_1 _14168_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._88_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._01_ ));
 sky130_fd_sc_hd__dfxtp_1 _14169_ (.CLK(clknet_leaf_132_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14170_ (.CLK(clknet_leaf_132_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14171_ (.CLK(clknet_leaf_132_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14172_ (.CLK(clknet_leaf_133_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14173_ (.CLK(clknet_leaf_132_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14174_ (.CLK(clknet_leaf_133_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14175_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14176_ (.CLK(clknet_leaf_132_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14177_ (.CLK(clknet_leaf_132_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14178_ (.CLK(clknet_leaf_132_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14179_ (.CLK(clknet_leaf_131_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14180_ (.CLK(clknet_leaf_120_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14181_ (.CLK(clknet_leaf_132_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14182_ (.CLK(clknet_leaf_132_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14183_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14184_ (.CLK(clknet_leaf_132_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14185_ (.CLK(clknet_leaf_133_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14186_ (.CLK(clknet_leaf_133_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14187_ (.CLK(clknet_leaf_133_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14188_ (.CLK(clknet_leaf_133_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14189_ (.CLK(clknet_leaf_133_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14190_ (.CLK(clknet_leaf_143_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14191_ (.CLK(clknet_leaf_143_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._35_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._02_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14192_ (.CLK(clknet_leaf_145_clk),
    .D(_00353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._24_ ));
 sky130_fd_sc_hd__dfxtp_2 _14193_ (.CLK(clknet_leaf_143_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._42_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._06_ ));
 sky130_fd_sc_hd__dfxtp_1 _14194_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._07_ ));
 sky130_fd_sc_hd__dfxtp_1 _14195_ (.CLK(clknet_leaf_132_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._48_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._08_ ));
 sky130_fd_sc_hd__dfxtp_1 _14196_ (.CLK(clknet_leaf_132_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._50_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._09_ ));
 sky130_fd_sc_hd__dfxtp_1 _14197_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._56_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i._31_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14198_ (.CLK(clknet_leaf_134_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14199_ (.CLK(clknet_leaf_134_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14200_ (.CLK(clknet_leaf_134_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14201_ (.CLK(clknet_leaf_133_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14202_ (.CLK(clknet_leaf_134_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14203_ (.CLK(clknet_leaf_134_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14204_ (.CLK(clknet_leaf_141_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14205_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14206_ (.CLK(clknet_leaf_141_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14207_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._59_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._12_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14208_ (.CLK(clknet_leaf_141_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._67_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._13_ ));
 sky130_fd_sc_hd__dfxtp_1 _14209_ (.CLK(clknet_leaf_142_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._69_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._14_ ));
 sky130_fd_sc_hd__dfxtp_1 _14210_ (.CLK(clknet_leaf_134_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._74_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.lzoc_inst._15_ ));
 sky130_fd_sc_hd__dfxtp_1 _14211_ (.CLK(clknet_leaf_89_clk),
    .D(\sa_inst.sak._19_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14212_ (.CLK(clknet_leaf_89_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w2_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14213_ (.CLK(clknet_leaf_88_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w3_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14214_ (.CLK(clknet_leaf_88_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w4_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14215_ (.CLK(clknet_leaf_88_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w5_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14216_ (.CLK(clknet_leaf_88_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w6_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14217_ (.CLK(clknet_leaf_88_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w7_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14218_ (.CLK(clknet_leaf_88_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w8_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14219_ (.CLK(clknet_leaf_88_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w9_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14220_ (.CLK(clknet_leaf_88_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w10_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14221_ (.CLK(clknet_leaf_182_clk),
    .D(_00354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14222_ (.CLK(clknet_leaf_187_clk),
    .D(_00355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14223_ (.CLK(clknet_leaf_180_clk),
    .D(_00356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14224_ (.CLK(clknet_leaf_180_clk),
    .D(_00357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14225_ (.CLK(clknet_leaf_180_clk),
    .D(_00358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14226_ (.CLK(clknet_leaf_173_clk),
    .D(_00359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14227_ (.CLK(clknet_leaf_173_clk),
    .D(_00360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14228_ (.CLK(clknet_leaf_153_clk),
    .D(_00361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14229_ (.CLK(clknet_leaf_174_clk),
    .D(_00362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14230_ (.CLK(clknet_leaf_153_clk),
    .D(_00363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14231_ (.CLK(clknet_leaf_151_clk),
    .D(_00364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14232_ (.CLK(clknet_leaf_151_clk),
    .D(_00365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14233_ (.CLK(clknet_leaf_151_clk),
    .D(_00366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14234_ (.CLK(clknet_leaf_177_clk),
    .D(_00367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14235_ (.CLK(clknet_leaf_177_clk),
    .D(_00368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14236_ (.CLK(clknet_leaf_3_clk),
    .D(_00369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14237_ (.CLK(clknet_leaf_3_clk),
    .D(_00370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14238_ (.CLK(clknet_leaf_0_clk),
    .D(_00371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14239_ (.CLK(clknet_leaf_0_clk),
    .D(_00372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14240_ (.CLK(clknet_leaf_0_clk),
    .D(_00373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14241_ (.CLK(clknet_leaf_191_clk),
    .D(_00374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14242_ (.CLK(clknet_leaf_191_clk),
    .D(_00375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14243_ (.CLK(clknet_leaf_189_clk),
    .D(_00376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14244_ (.CLK(clknet_leaf_189_clk),
    .D(_00377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14245_ (.CLK(clknet_leaf_86_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14246_ (.CLK(clknet_leaf_86_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14247_ (.CLK(clknet_leaf_92_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14248_ (.CLK(clknet_leaf_92_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14249_ (.CLK(clknet_leaf_91_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14250_ (.CLK(clknet_leaf_92_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14251_ (.CLK(clknet_leaf_91_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14252_ (.CLK(clknet_leaf_86_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14253_ (.CLK(clknet_leaf_86_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14254_ (.CLK(clknet_leaf_86_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14255_ (.CLK(clknet_leaf_86_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14256_ (.CLK(clknet_leaf_86_clk),
    .D(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._3_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:2.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14257_ (.CLK(clknet_leaf_181_clk),
    .D(_00378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14258_ (.CLK(clknet_leaf_187_clk),
    .D(_00379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14259_ (.CLK(clknet_leaf_178_clk),
    .D(_00380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14260_ (.CLK(clknet_leaf_178_clk),
    .D(_00381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14261_ (.CLK(clknet_leaf_178_clk),
    .D(_00382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14262_ (.CLK(clknet_leaf_159_clk),
    .D(_00383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14263_ (.CLK(clknet_leaf_154_clk),
    .D(_00384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14264_ (.CLK(clknet_leaf_157_clk),
    .D(_00385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14265_ (.CLK(clknet_leaf_157_clk),
    .D(_00386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14266_ (.CLK(clknet_leaf_156_clk),
    .D(_00387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14267_ (.CLK(clknet_leaf_149_clk),
    .D(_00388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14268_ (.CLK(clknet_leaf_148_clk),
    .D(_00389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14269_ (.CLK(clknet_leaf_147_clk),
    .D(_00390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14270_ (.CLK(clknet_leaf_147_clk),
    .D(_00391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14271_ (.CLK(clknet_leaf_147_clk),
    .D(_00392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14272_ (.CLK(clknet_leaf_4_clk),
    .D(_00393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14273_ (.CLK(clknet_leaf_4_clk),
    .D(_00394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14274_ (.CLK(clknet_leaf_5_clk),
    .D(_00395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14275_ (.CLK(clknet_leaf_5_clk),
    .D(_00396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14276_ (.CLK(clknet_leaf_3_clk),
    .D(_00397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14277_ (.CLK(clknet_leaf_190_clk),
    .D(_00398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14278_ (.CLK(clknet_leaf_190_clk),
    .D(_00399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14279_ (.CLK(clknet_leaf_188_clk),
    .D(_00400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14280_ (.CLK(clknet_leaf_188_clk),
    .D(_00401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14281_ (.CLK(clknet_leaf_138_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.rshift._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.rshift._11_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14282_ (.CLK(clknet_leaf_137_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._35_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.rshift._22_ ));
 sky130_fd_sc_hd__dfxtp_1 _14283_ (.CLK(clknet_leaf_137_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.rshift._04_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.rshift._25_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14284_ (.CLK(clknet_leaf_137_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.rshift._04_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.rshift._25_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14285_ (.CLK(clknet_leaf_137_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.rshift._04_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.rshift._25_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14286_ (.CLK(clknet_leaf_137_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.rshift._04_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.rshift._25_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14287_ (.CLK(clknet_leaf_138_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.rshift._10_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.rshift._26_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14288_ (.CLK(clknet_leaf_138_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.rshift._10_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.rshift._26_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14289_ (.CLK(clknet_leaf_137_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.rshift._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.rshift._27_ ));
 sky130_fd_sc_hd__dfxtp_1 _14290_ (.CLK(clknet_leaf_138_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.rshift._17_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.rshift._28_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14291_ (.CLK(clknet_leaf_138_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i.rshift._28_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.rshift._18_ ));
 sky130_fd_sc_hd__dfxtp_1 _14292_ (.CLK(clknet_leaf_138_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._35_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.rshift._00_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14293_ (.CLK(clknet_leaf_137_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._35_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.rshift._00_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14294_ (.CLK(clknet_leaf_137_clk),
    .D(\sa_inst.cols_l2a:2.l2a_i._35_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:2.l2a_i.rshift._00_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14295_ (.CLK(clknet_leaf_183_clk),
    .D(_00402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14296_ (.CLK(clknet_leaf_182_clk),
    .D(_00403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14297_ (.CLK(clknet_leaf_183_clk),
    .D(_00404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14298_ (.CLK(clknet_leaf_176_clk),
    .D(_00405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14299_ (.CLK(clknet_leaf_179_clk),
    .D(_00406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14300_ (.CLK(clknet_leaf_153_clk),
    .D(_00407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14301_ (.CLK(clknet_leaf_175_clk),
    .D(_00408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14302_ (.CLK(clknet_leaf_153_clk),
    .D(_00409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14303_ (.CLK(clknet_leaf_153_clk),
    .D(_00410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14304_ (.CLK(clknet_leaf_153_clk),
    .D(_00411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14305_ (.CLK(clknet_leaf_152_clk),
    .D(_00412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14306_ (.CLK(clknet_leaf_151_clk),
    .D(_00413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14307_ (.CLK(clknet_leaf_152_clk),
    .D(_00414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14308_ (.CLK(clknet_leaf_151_clk),
    .D(_00415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14309_ (.CLK(clknet_leaf_151_clk),
    .D(_00416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14310_ (.CLK(clknet_leaf_3_clk),
    .D(_00417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14311_ (.CLK(clknet_leaf_185_clk),
    .D(_00418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14312_ (.CLK(clknet_leaf_0_clk),
    .D(_00419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14313_ (.CLK(clknet_leaf_0_clk),
    .D(_00420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14314_ (.CLK(clknet_leaf_0_clk),
    .D(_00421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14315_ (.CLK(clknet_leaf_191_clk),
    .D(_00422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14316_ (.CLK(clknet_leaf_191_clk),
    .D(_00423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14317_ (.CLK(clknet_leaf_186_clk),
    .D(_00424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14318_ (.CLK(clknet_leaf_189_clk),
    .D(_00425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[8][23] ));
 sky130_fd_sc_hd__dfxtp_2 _14319_ (.CLK(clknet_leaf_13_clk),
    .D(\sa_inst._12_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._00_ ));
 sky130_fd_sc_hd__dfxtp_1 _14320_ (.CLK(clknet_leaf_166_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._26_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._27_ ));
 sky130_fd_sc_hd__dfxtp_1 _14321_ (.CLK(clknet_leaf_167_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._25_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._26_ ));
 sky130_fd_sc_hd__dfxtp_1 _14322_ (.CLK(clknet_leaf_168_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._24_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._25_ ));
 sky130_fd_sc_hd__dfxtp_1 _14323_ (.CLK(clknet_leaf_79_clk),
    .D(_00426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14324_ (.CLK(clknet_leaf_79_clk),
    .D(_00427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14325_ (.CLK(clknet_leaf_79_clk),
    .D(_00428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14326_ (.CLK(clknet_leaf_79_clk),
    .D(_00429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._09_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14327_ (.CLK(clknet_leaf_158_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._21_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._23_ ));
 sky130_fd_sc_hd__dfxtp_1 _14328_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._20_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._21_ ));
 sky130_fd_sc_hd__dfxtp_1 _14329_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._19_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._20_ ));
 sky130_fd_sc_hd__dfxtp_1 _14330_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._18_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._19_ ));
 sky130_fd_sc_hd__dfxtp_1 _14331_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._17_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._18_ ));
 sky130_fd_sc_hd__dfxtp_1 _14332_ (.CLK(clknet_leaf_162_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._16_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._17_ ));
 sky130_fd_sc_hd__dfxtp_1 _14333_ (.CLK(clknet_leaf_162_clk),
    .D(\sa_inst._12_[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._16_ ));
 sky130_fd_sc_hd__dfxtp_1 _14334_ (.CLK(clknet_leaf_160_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._46_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._15_ ));
 sky130_fd_sc_hd__dfxtp_1 _14335_ (.CLK(clknet_leaf_165_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._13_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._14_ ));
 sky130_fd_sc_hd__dfxtp_1 _14336_ (.CLK(clknet_leaf_165_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._40_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._13_ ));
 sky130_fd_sc_hd__dfxtp_1 _14337_ (.CLK(clknet_leaf_160_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._08_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._09_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14338_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._08_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._09_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14339_ (.CLK(clknet_leaf_160_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._08_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._09_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14340_ (.CLK(clknet_leaf_160_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._08_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._09_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14341_ (.CLK(clknet_leaf_160_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._08_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._09_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14342_ (.CLK(clknet_leaf_160_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._08_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._09_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14343_ (.CLK(clknet_leaf_160_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._08_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._09_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14344_ (.CLK(clknet_leaf_166_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._07_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._08_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14345_ (.CLK(clknet_leaf_160_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._07_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._08_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14346_ (.CLK(clknet_leaf_166_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._07_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._08_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14347_ (.CLK(clknet_leaf_166_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._07_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._08_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14348_ (.CLK(clknet_leaf_166_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._07_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._08_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14349_ (.CLK(clknet_leaf_166_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._07_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._08_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14350_ (.CLK(clknet_leaf_160_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._07_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._08_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14351_ (.CLK(clknet_leaf_165_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._40_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._07_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14352_ (.CLK(clknet_leaf_166_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._40_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._07_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14353_ (.CLK(clknet_leaf_166_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._40_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._07_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14354_ (.CLK(clknet_leaf_166_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._40_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._07_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14355_ (.CLK(clknet_leaf_166_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._40_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._07_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14356_ (.CLK(clknet_leaf_166_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._40_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._07_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14357_ (.CLK(clknet_leaf_166_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._37_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._07_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14358_ (.CLK(clknet_leaf_168_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._31_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._06_ ));
 sky130_fd_sc_hd__dfxtp_1 _14359_ (.CLK(clknet_leaf_167_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._31_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._05_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14360_ (.CLK(clknet_leaf_167_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._31_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._05_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14361_ (.CLK(clknet_leaf_168_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._31_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._05_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14362_ (.CLK(clknet_leaf_168_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._31_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._05_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14363_ (.CLK(clknet_leaf_165_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._03_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._04_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14364_ (.CLK(clknet_leaf_165_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._02_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._03_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14365_ (.CLK(clknet_leaf_168_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._29_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._02_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14366_ (.CLK(clknet_leaf_168_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._29_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._02_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14367_ (.CLK(clknet_leaf_168_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._29_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._02_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14368_ (.CLK(clknet_leaf_168_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._29_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._02_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14369_ (.CLK(clknet_leaf_168_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._29_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._02_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14370_ (.CLK(clknet_leaf_168_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._29_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._02_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14371_ (.CLK(clknet_leaf_167_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._57_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._01_ ));
 sky130_fd_sc_hd__dfxtp_1 _14372_ (.CLK(clknet_leaf_167_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._56_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._57_ ));
 sky130_fd_sc_hd__dfxtp_1 _14373_ (.CLK(clknet_leaf_167_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._30_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._56_ ));
 sky130_fd_sc_hd__dfxtp_1 _14374_ (.CLK(clknet_leaf_159_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._54_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._55_ ));
 sky130_fd_sc_hd__dfxtp_1 _14375_ (.CLK(clknet_leaf_167_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._44_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._54_ ));
 sky130_fd_sc_hd__dfxtp_1 _14376_ (.CLK(clknet_leaf_167_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._33_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._44_ ));
 sky130_fd_sc_hd__dfxtp_1 _14377_ (.CLK(clknet_leaf_167_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._22_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._33_ ));
 sky130_fd_sc_hd__dfxtp_1 _14378_ (.CLK(clknet_leaf_170_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._11_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._22_ ));
 sky130_fd_sc_hd__dfxtp_1 _14379_ (.CLK(clknet_leaf_170_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._00_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._11_ ));
 sky130_fd_sc_hd__dfxtp_1 _14380_ (.CLK(clknet_leaf_17_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._23_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._33_ ));
 sky130_fd_sc_hd__dfxtp_1 _14381_ (.CLK(clknet_leaf_17_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._33_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._44_ ));
 sky130_fd_sc_hd__dfxtp_1 _14382_ (.CLK(clknet_leaf_17_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._44_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._55_ ));
 sky130_fd_sc_hd__dfxtp_1 _14383_ (.CLK(clknet_leaf_16_clk),
    .D(_00430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._05_ ));
 sky130_fd_sc_hd__dfxtp_1 _14384_ (.CLK(clknet_leaf_17_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._31_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._88_ ));
 sky130_fd_sc_hd__dfxtp_1 _14385_ (.CLK(clknet_leaf_16_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._88_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._01_ ));
 sky130_fd_sc_hd__dfxtp_1 _14386_ (.CLK(clknet_leaf_16_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14387_ (.CLK(clknet_leaf_16_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14388_ (.CLK(clknet_leaf_16_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14389_ (.CLK(clknet_leaf_16_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14390_ (.CLK(clknet_leaf_15_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14391_ (.CLK(clknet_leaf_170_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14392_ (.CLK(clknet_leaf_15_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14393_ (.CLK(clknet_leaf_15_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14394_ (.CLK(clknet_leaf_16_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14395_ (.CLK(clknet_leaf_16_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14396_ (.CLK(clknet_leaf_16_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14397_ (.CLK(clknet_leaf_17_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14398_ (.CLK(clknet_leaf_15_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14399_ (.CLK(clknet_leaf_170_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14400_ (.CLK(clknet_leaf_15_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14401_ (.CLK(clknet_leaf_15_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14402_ (.CLK(clknet_leaf_15_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14403_ (.CLK(clknet_leaf_15_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14404_ (.CLK(clknet_leaf_15_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14405_ (.CLK(clknet_leaf_15_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14406_ (.CLK(clknet_leaf_15_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14407_ (.CLK(clknet_leaf_15_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14408_ (.CLK(clknet_leaf_15_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._35_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._02_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14409_ (.CLK(clknet_leaf_168_clk),
    .D(_00431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._24_ ));
 sky130_fd_sc_hd__dfxtp_2 _14410_ (.CLK(clknet_leaf_15_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._42_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._06_ ));
 sky130_fd_sc_hd__dfxtp_1 _14411_ (.CLK(clknet_leaf_16_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._06_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._07_ ));
 sky130_fd_sc_hd__dfxtp_1 _14412_ (.CLK(clknet_leaf_16_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._48_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._08_ ));
 sky130_fd_sc_hd__dfxtp_1 _14413_ (.CLK(clknet_leaf_16_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._50_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._09_ ));
 sky130_fd_sc_hd__dfxtp_1 _14414_ (.CLK(clknet_leaf_169_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._56_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i._31_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14415_ (.CLK(clknet_leaf_169_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14416_ (.CLK(clknet_leaf_169_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14417_ (.CLK(clknet_leaf_170_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14418_ (.CLK(clknet_leaf_168_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14419_ (.CLK(clknet_leaf_170_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14420_ (.CLK(clknet_leaf_170_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14421_ (.CLK(clknet_leaf_169_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14422_ (.CLK(clknet_leaf_169_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14423_ (.CLK(clknet_leaf_170_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14424_ (.CLK(clknet_leaf_169_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._59_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._12_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14425_ (.CLK(clknet_leaf_168_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._67_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._13_ ));
 sky130_fd_sc_hd__dfxtp_1 _14426_ (.CLK(clknet_leaf_170_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._69_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._14_ ));
 sky130_fd_sc_hd__dfxtp_1 _14427_ (.CLK(clknet_leaf_167_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._74_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.lzoc_inst._15_ ));
 sky130_fd_sc_hd__dfxtp_1 _14428_ (.CLK(clknet_leaf_55_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._14_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14429_ (.CLK(clknet_leaf_54_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._14_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14430_ (.CLK(clknet_leaf_46_clk),
    .D(\sa_inst._05_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak._00_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14431_ (.CLK(clknet_leaf_44_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w2_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14432_ (.CLK(clknet_leaf_47_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w3_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14433_ (.CLK(clknet_leaf_44_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w4_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14434_ (.CLK(clknet_leaf_45_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w5_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14435_ (.CLK(clknet_leaf_44_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w6_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14436_ (.CLK(clknet_leaf_45_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w7_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14437_ (.CLK(clknet_leaf_45_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w8_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14438_ (.CLK(clknet_leaf_45_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w9_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14439_ (.CLK(clknet_leaf_45_clk),
    .D(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_inst.bh33_w10_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:1.cols:1.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14440_ (.CLK(clknet_leaf_88_clk),
    .D(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_inst.bh33_w11_0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.sak.rows:3.cols:3.pe_ij.s3fdp_inst.significand_product_shifter_inst._1_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14441_ (.CLK(clknet_leaf_183_clk),
    .D(_00432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14442_ (.CLK(clknet_leaf_187_clk),
    .D(_00433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14443_ (.CLK(clknet_leaf_176_clk),
    .D(_00434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14444_ (.CLK(clknet_leaf_177_clk),
    .D(_00435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14445_ (.CLK(clknet_leaf_176_clk),
    .D(_00436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14446_ (.CLK(clknet_leaf_153_clk),
    .D(_00437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14447_ (.CLK(clknet_leaf_153_clk),
    .D(_00438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14448_ (.CLK(clknet_leaf_155_clk),
    .D(_00439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14449_ (.CLK(clknet_leaf_155_clk),
    .D(_00440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14450_ (.CLK(clknet_leaf_155_clk),
    .D(_00441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14451_ (.CLK(clknet_leaf_152_clk),
    .D(_00442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14452_ (.CLK(clknet_leaf_149_clk),
    .D(_00443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14453_ (.CLK(clknet_leaf_145_clk),
    .D(_00444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14454_ (.CLK(clknet_leaf_145_clk),
    .D(_00445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14455_ (.CLK(clknet_leaf_148_clk),
    .D(_00446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14456_ (.CLK(clknet_leaf_186_clk),
    .D(_00447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14457_ (.CLK(clknet_leaf_185_clk),
    .D(_00448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14458_ (.CLK(clknet_leaf_2_clk),
    .D(_00449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14459_ (.CLK(clknet_leaf_2_clk),
    .D(_00450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14460_ (.CLK(clknet_leaf_192_clk),
    .D(_00451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14461_ (.CLK(clknet_leaf_191_clk),
    .D(_00452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14462_ (.CLK(clknet_leaf_189_clk),
    .D(_00453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14463_ (.CLK(clknet_leaf_186_clk),
    .D(_00454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14464_ (.CLK(clknet_leaf_189_clk),
    .D(_00455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14465_ (.CLK(clknet_leaf_183_clk),
    .D(_00456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14466_ (.CLK(clknet_leaf_187_clk),
    .D(_00457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14467_ (.CLK(clknet_leaf_183_clk),
    .D(_00458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14468_ (.CLK(clknet_leaf_179_clk),
    .D(_00459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14469_ (.CLK(clknet_leaf_179_clk),
    .D(_00460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14470_ (.CLK(clknet_leaf_174_clk),
    .D(_00461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14471_ (.CLK(clknet_leaf_175_clk),
    .D(_00462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14472_ (.CLK(clknet_leaf_153_clk),
    .D(_00463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14473_ (.CLK(clknet_leaf_175_clk),
    .D(_00464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14474_ (.CLK(clknet_leaf_153_clk),
    .D(_00465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14475_ (.CLK(clknet_leaf_152_clk),
    .D(_00466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14476_ (.CLK(clknet_leaf_151_clk),
    .D(_00467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14477_ (.CLK(clknet_leaf_152_clk),
    .D(_00468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14478_ (.CLK(clknet_leaf_177_clk),
    .D(_00469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14479_ (.CLK(clknet_leaf_151_clk),
    .D(_00470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14480_ (.CLK(clknet_leaf_3_clk),
    .D(_00471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14481_ (.CLK(clknet_leaf_185_clk),
    .D(_00472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14482_ (.CLK(clknet_leaf_0_clk),
    .D(_00473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14483_ (.CLK(clknet_leaf_0_clk),
    .D(_00474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14484_ (.CLK(clknet_leaf_0_clk),
    .D(_00475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14485_ (.CLK(clknet_leaf_191_clk),
    .D(_00476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14486_ (.CLK(clknet_leaf_191_clk),
    .D(_00477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14487_ (.CLK(clknet_leaf_186_clk),
    .D(_00478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14488_ (.CLK(clknet_leaf_189_clk),
    .D(_00479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14489_ (.CLK(clknet_leaf_184_clk),
    .D(_00480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14490_ (.CLK(clknet_leaf_186_clk),
    .D(_00481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14491_ (.CLK(clknet_leaf_172_clk),
    .D(_00482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14492_ (.CLK(clknet_leaf_172_clk),
    .D(_00483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14493_ (.CLK(clknet_leaf_176_clk),
    .D(_00484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14494_ (.CLK(clknet_leaf_153_clk),
    .D(_00485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14495_ (.CLK(clknet_leaf_153_clk),
    .D(_00486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14496_ (.CLK(clknet_leaf_155_clk),
    .D(_00487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14497_ (.CLK(clknet_leaf_144_clk),
    .D(_00488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14498_ (.CLK(clknet_leaf_155_clk),
    .D(_00489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14499_ (.CLK(clknet_leaf_152_clk),
    .D(_00490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14500_ (.CLK(clknet_leaf_152_clk),
    .D(_00491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14501_ (.CLK(clknet_leaf_145_clk),
    .D(_00492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14502_ (.CLK(clknet_leaf_145_clk),
    .D(_00493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14503_ (.CLK(clknet_leaf_145_clk),
    .D(_00494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14504_ (.CLK(clknet_leaf_2_clk),
    .D(_00495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14505_ (.CLK(clknet_leaf_186_clk),
    .D(_00496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14506_ (.CLK(clknet_leaf_2_clk),
    .D(_00497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14507_ (.CLK(clknet_leaf_192_clk),
    .D(_00498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14508_ (.CLK(clknet_leaf_192_clk),
    .D(_00499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14509_ (.CLK(clknet_leaf_191_clk),
    .D(_00500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14510_ (.CLK(clknet_leaf_0_clk),
    .D(_00501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14511_ (.CLK(clknet_leaf_186_clk),
    .D(_00502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14512_ (.CLK(clknet_leaf_2_clk),
    .D(_00503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[6][23] ));
 sky130_fd_sc_hd__dfxtp_2 _14513_ (.CLK(clknet_leaf_146_clk),
    .D(_00504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.WR_DATA[8] ));
 sky130_fd_sc_hd__dfxtp_2 _14514_ (.CLK(clknet_leaf_146_clk),
    .D(_00505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.WR_DATA[9] ));
 sky130_fd_sc_hd__dfxtp_2 _14515_ (.CLK(clknet_leaf_146_clk),
    .D(_00506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.WR_DATA[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14516_ (.CLK(clknet_leaf_146_clk),
    .D(_00507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.WR_DATA[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14517_ (.CLK(clknet_leaf_146_clk),
    .D(_00508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.WR_DATA[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14518_ (.CLK(clknet_leaf_147_clk),
    .D(_00509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.WR_DATA[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14519_ (.CLK(clknet_leaf_146_clk),
    .D(_00510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.WR_DATA[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14520_ (.CLK(clknet_leaf_163_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.rshift._00_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.rshift._11_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14521_ (.CLK(clknet_leaf_165_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._35_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.rshift._22_ ));
 sky130_fd_sc_hd__dfxtp_1 _14522_ (.CLK(clknet_leaf_164_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.rshift._04_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.rshift._25_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14523_ (.CLK(clknet_leaf_165_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.rshift._04_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.rshift._25_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14524_ (.CLK(clknet_leaf_165_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.rshift._04_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.rshift._25_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14525_ (.CLK(clknet_leaf_165_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.rshift._04_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.rshift._25_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14526_ (.CLK(clknet_leaf_164_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.rshift._10_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.rshift._26_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14527_ (.CLK(clknet_leaf_164_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.rshift._10_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.rshift._26_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14528_ (.CLK(clknet_leaf_165_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.rshift._14_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.rshift._27_ ));
 sky130_fd_sc_hd__dfxtp_1 _14529_ (.CLK(clknet_leaf_164_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.rshift._17_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.rshift._28_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14530_ (.CLK(clknet_leaf_163_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i.rshift._28_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.rshift._18_ ));
 sky130_fd_sc_hd__dfxtp_1 _14531_ (.CLK(clknet_leaf_181_clk),
    .D(_00511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14532_ (.CLK(clknet_leaf_188_clk),
    .D(_00512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14533_ (.CLK(clknet_leaf_181_clk),
    .D(_00513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14534_ (.CLK(clknet_leaf_180_clk),
    .D(_00514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14535_ (.CLK(clknet_leaf_180_clk),
    .D(_00515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14536_ (.CLK(clknet_leaf_167_clk),
    .D(_00516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14537_ (.CLK(clknet_leaf_173_clk),
    .D(_00517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14538_ (.CLK(clknet_leaf_160_clk),
    .D(_00518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14539_ (.CLK(clknet_leaf_174_clk),
    .D(_00519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14540_ (.CLK(clknet_leaf_154_clk),
    .D(_00520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14541_ (.CLK(clknet_leaf_150_clk),
    .D(_00521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14542_ (.CLK(clknet_leaf_151_clk),
    .D(_00522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14543_ (.CLK(clknet_leaf_151_clk),
    .D(_00523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14544_ (.CLK(clknet_leaf_178_clk),
    .D(_00524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14545_ (.CLK(clknet_leaf_177_clk),
    .D(_00525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14546_ (.CLK(clknet_leaf_4_clk),
    .D(_00526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14547_ (.CLK(clknet_leaf_4_clk),
    .D(_00527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14548_ (.CLK(clknet_leaf_6_clk),
    .D(_00528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14549_ (.CLK(clknet_leaf_6_clk),
    .D(_00529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14550_ (.CLK(clknet_leaf_1_clk),
    .D(_00530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14551_ (.CLK(clknet_leaf_190_clk),
    .D(_00531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14552_ (.CLK(clknet_leaf_190_clk),
    .D(_00532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14553_ (.CLK(clknet_leaf_188_clk),
    .D(_00533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14554_ (.CLK(clknet_leaf_188_clk),
    .D(_00534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14555_ (.CLK(clknet_leaf_164_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._35_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.rshift._00_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14556_ (.CLK(clknet_leaf_165_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._35_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.rshift._00_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14557_ (.CLK(clknet_leaf_165_clk),
    .D(\sa_inst.cols_l2a:1.l2a_i._35_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_l2a:1.l2a_i.rshift._00_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14558_ (.CLK(clknet_leaf_184_clk),
    .D(_00535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14559_ (.CLK(clknet_leaf_184_clk),
    .D(_00536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14560_ (.CLK(clknet_leaf_176_clk),
    .D(_00537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14561_ (.CLK(clknet_leaf_177_clk),
    .D(_00538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14562_ (.CLK(clknet_leaf_175_clk),
    .D(_00539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14563_ (.CLK(clknet_leaf_155_clk),
    .D(_00540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14564_ (.CLK(clknet_leaf_152_clk),
    .D(_00541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14565_ (.CLK(clknet_leaf_144_clk),
    .D(_00542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14566_ (.CLK(clknet_leaf_144_clk),
    .D(_00543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14567_ (.CLK(clknet_leaf_155_clk),
    .D(_00544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14568_ (.CLK(clknet_leaf_152_clk),
    .D(_00545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14569_ (.CLK(clknet_leaf_149_clk),
    .D(_00546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14570_ (.CLK(clknet_leaf_145_clk),
    .D(_00547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14571_ (.CLK(clknet_leaf_144_clk),
    .D(_00548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14572_ (.CLK(clknet_leaf_145_clk),
    .D(_00549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14573_ (.CLK(clknet_leaf_186_clk),
    .D(_00550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14574_ (.CLK(clknet_leaf_185_clk),
    .D(_00551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14575_ (.CLK(clknet_leaf_2_clk),
    .D(_00552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14576_ (.CLK(clknet_leaf_2_clk),
    .D(_00553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14577_ (.CLK(clknet_leaf_192_clk),
    .D(_00554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14578_ (.CLK(clknet_leaf_192_clk),
    .D(_00555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14579_ (.CLK(clknet_leaf_192_clk),
    .D(_00556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14580_ (.CLK(clknet_leaf_186_clk),
    .D(_00557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14581_ (.CLK(clknet_leaf_186_clk),
    .D(_00558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14582_ (.CLK(clknet_leaf_80_clk),
    .D(\sa_inst._17_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:3.a2s3_j._00_ ));
 sky130_fd_sc_hd__dfxtp_1 _14583_ (.CLK(clknet_leaf_80_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j.43$func$/openlane/designs/teras/src/arith_to_s3.v:95$95.$result[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:3.a2s3_j._15_[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14584_ (.CLK(clknet_leaf_79_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j._19_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._07_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14585_ (.CLK(clknet_leaf_79_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j._07_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:3.a2s3_j._19_ ));
 sky130_fd_sc_hd__dfxtp_2 _14586_ (.CLK(clknet_leaf_79_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j._17_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._07_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14587_ (.CLK(clknet_leaf_79_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:3.a2s3_j._17_ ));
 sky130_fd_sc_hd__dfxtp_2 _14588_ (.CLK(clknet_leaf_83_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j._00_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._07_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14589_ (.CLK(clknet_leaf_81_clk),
    .D(\sa_inst._17_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._00_ ));
 sky130_fd_sc_hd__dfxtp_1 _14590_ (.CLK(clknet_leaf_79_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._11_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._08_ ));
 sky130_fd_sc_hd__dfxtp_1 _14591_ (.CLK(clknet_leaf_55_clk),
    .D(_00559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14592_ (.CLK(clknet_leaf_55_clk),
    .D(_00560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14593_ (.CLK(clknet_leaf_55_clk),
    .D(_00561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14594_ (.CLK(clknet_leaf_54_clk),
    .D(_00562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._09_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14595_ (.CLK(clknet_leaf_80_clk),
    .D(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._01_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:3.a2s3_j.lzoc._10_ ));
 sky130_fd_sc_hd__dfxtp_1 _14596_ (.CLK(clknet_leaf_184_clk),
    .D(_00563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14597_ (.CLK(clknet_leaf_184_clk),
    .D(_00564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14598_ (.CLK(clknet_leaf_176_clk),
    .D(_00565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14599_ (.CLK(clknet_leaf_175_clk),
    .D(_00566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14600_ (.CLK(clknet_leaf_175_clk),
    .D(_00567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14601_ (.CLK(clknet_leaf_155_clk),
    .D(_00568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14602_ (.CLK(clknet_leaf_152_clk),
    .D(_00569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14603_ (.CLK(clknet_leaf_144_clk),
    .D(_00570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14604_ (.CLK(clknet_leaf_144_clk),
    .D(_00571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14605_ (.CLK(clknet_leaf_144_clk),
    .D(_00572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14606_ (.CLK(clknet_leaf_149_clk),
    .D(_00573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14607_ (.CLK(clknet_leaf_148_clk),
    .D(_00574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14608_ (.CLK(clknet_leaf_146_clk),
    .D(_00575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14609_ (.CLK(clknet_leaf_145_clk),
    .D(_00576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14610_ (.CLK(clknet_leaf_145_clk),
    .D(_00577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14611_ (.CLK(clknet_leaf_186_clk),
    .D(_00578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14612_ (.CLK(clknet_leaf_185_clk),
    .D(_00579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14613_ (.CLK(clknet_leaf_2_clk),
    .D(_00580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14614_ (.CLK(clknet_leaf_2_clk),
    .D(_00581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14615_ (.CLK(clknet_leaf_2_clk),
    .D(_00582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14616_ (.CLK(clknet_leaf_191_clk),
    .D(_00583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14617_ (.CLK(clknet_leaf_191_clk),
    .D(_00584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14618_ (.CLK(clknet_leaf_186_clk),
    .D(_00585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14619_ (.CLK(clknet_leaf_186_clk),
    .D(_00586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14620_ (.CLK(clknet_leaf_78_clk),
    .D(\sa_inst._00_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:2.a2s3_j._00_ ));
 sky130_fd_sc_hd__dfxtp_4 _14621_ (.CLK(clknet_leaf_56_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j._15_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._06_[0] ));
 sky130_fd_sc_hd__dfxtp_2 _14622_ (.CLK(clknet_leaf_56_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j._15_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:2.a2s3_j._23_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14623_ (.CLK(clknet_leaf_61_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j._15_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:2.a2s3_j._23_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14624_ (.CLK(clknet_leaf_61_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j._15_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:2.a2s3_j._23_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14625_ (.CLK(clknet_leaf_53_clk),
    .D(_00587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14626_ (.CLK(clknet_leaf_52_clk),
    .D(_00588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14627_ (.CLK(clknet_leaf_52_clk),
    .D(_00589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14628_ (.CLK(clknet_leaf_51_clk),
    .D(_00590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._09_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14629_ (.CLK(clknet_leaf_56_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j.43$func$/openlane/designs/teras/src/arith_to_s3.v:95$95.$result[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:2.a2s3_j._15_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14630_ (.CLK(clknet_leaf_55_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j._19_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._06_[9] ));
 sky130_fd_sc_hd__dfxtp_2 _14631_ (.CLK(clknet_leaf_78_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j._00_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._06_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14632_ (.CLK(clknet_leaf_55_clk),
    .D(\sa_inst._00_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._00_ ));
 sky130_fd_sc_hd__dfxtp_1 _14633_ (.CLK(clknet_leaf_53_clk),
    .D(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._11_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:2.a2s3_j.lzoc._08_ ));
 sky130_fd_sc_hd__dfxtp_2 _14634_ (.CLK(clknet_leaf_57_clk),
    .D(_00591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._06_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14635_ (.CLK(clknet_leaf_61_clk),
    .D(\sa_inst.arith_in_col_0[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:1.a2s3_j._00_ ));
 sky130_fd_sc_hd__dfxtp_1 _14636_ (.CLK(clknet_leaf_61_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j._00_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._05_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14637_ (.CLK(clknet_leaf_51_clk),
    .D(\sa_inst.arith_in_col_0[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._00_ ));
 sky130_fd_sc_hd__dfxtp_1 _14638_ (.CLK(clknet_leaf_52_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._11_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._08_ ));
 sky130_fd_sc_hd__dfxtp_1 _14639_ (.CLK(clknet_leaf_54_clk),
    .D(_00592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._00_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14640_ (.CLK(clknet_leaf_55_clk),
    .D(_00593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._00_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14641_ (.CLK(clknet_leaf_54_clk),
    .D(_00594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._00_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14642_ (.CLK(clknet_leaf_54_clk),
    .D(_00595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._00_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14643_ (.CLK(clknet_leaf_54_clk),
    .D(_00596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._00_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14644_ (.CLK(clknet_leaf_55_clk),
    .D(_00597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._00_[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14645_ (.CLK(clknet_leaf_56_clk),
    .D(_00598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._00_[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14646_ (.CLK(clknet_leaf_78_clk),
    .D(_00599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._00_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14647_ (.CLK(clknet_leaf_52_clk),
    .D(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._01_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst.cols_a2s3:1.a2s3_j.lzoc._10_ ));
 sky130_fd_sc_hd__dfxtp_1 _14648_ (.CLK(clknet_leaf_182_clk),
    .D(_00600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14649_ (.CLK(clknet_leaf_182_clk),
    .D(_00601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14650_ (.CLK(clknet_leaf_179_clk),
    .D(_00602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14651_ (.CLK(clknet_leaf_177_clk),
    .D(_00603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14652_ (.CLK(clknet_leaf_177_clk),
    .D(_00604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14653_ (.CLK(clknet_leaf_159_clk),
    .D(_00605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14654_ (.CLK(clknet_leaf_154_clk),
    .D(_00606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14655_ (.CLK(clknet_leaf_159_clk),
    .D(_00607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14656_ (.CLK(clknet_leaf_157_clk),
    .D(_00608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14657_ (.CLK(clknet_leaf_156_clk),
    .D(_00609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14658_ (.CLK(clknet_leaf_149_clk),
    .D(_00610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14659_ (.CLK(clknet_leaf_149_clk),
    .D(_00611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14660_ (.CLK(clknet_leaf_147_clk),
    .D(_00612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14661_ (.CLK(clknet_leaf_147_clk),
    .D(_00613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14662_ (.CLK(clknet_leaf_148_clk),
    .D(_00614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14663_ (.CLK(clknet_leaf_3_clk),
    .D(_00615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14664_ (.CLK(clknet_leaf_185_clk),
    .D(_00616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14665_ (.CLK(clknet_leaf_4_clk),
    .D(_00617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14666_ (.CLK(clknet_leaf_3_clk),
    .D(_00618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14667_ (.CLK(clknet_leaf_3_clk),
    .D(_00619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14668_ (.CLK(clknet_leaf_189_clk),
    .D(_00620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14669_ (.CLK(clknet_leaf_190_clk),
    .D(_00621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14670_ (.CLK(clknet_leaf_187_clk),
    .D(_00622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14671_ (.CLK(clknet_leaf_189_clk),
    .D(_00623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14672_ (.CLK(clknet_leaf_79_clk),
    .D(_00624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._11_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14673_ (.CLK(clknet_leaf_79_clk),
    .D(_00625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._11_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14674_ (.CLK(clknet_leaf_82_clk),
    .D(_00626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._11_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14675_ (.CLK(clknet_leaf_79_clk),
    .D(_00627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._11_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14676_ (.CLK(clknet_leaf_82_clk),
    .D(_00628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._11_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14677_ (.CLK(clknet_leaf_79_clk),
    .D(_00629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._11_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14678_ (.CLK(clknet_leaf_81_clk),
    .D(_00630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._11_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14679_ (.CLK(clknet_leaf_78_clk),
    .D(_00631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._11_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14680_ (.CLK(clknet_leaf_48_clk),
    .D(_00632_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._21_ ));
 sky130_fd_sc_hd__dfxtp_1 _14681_ (.CLK(clknet_leaf_79_clk),
    .D(\sa_inst._11_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._17_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14682_ (.CLK(clknet_leaf_79_clk),
    .D(\sa_inst._11_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._17_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14683_ (.CLK(clknet_leaf_82_clk),
    .D(\sa_inst._11_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._17_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14684_ (.CLK(clknet_leaf_79_clk),
    .D(\sa_inst._11_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._17_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14685_ (.CLK(clknet_leaf_82_clk),
    .D(\sa_inst._11_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._17_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14686_ (.CLK(clknet_leaf_79_clk),
    .D(\sa_inst._11_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._17_[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14687_ (.CLK(clknet_leaf_82_clk),
    .D(\sa_inst._11_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._17_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14688_ (.CLK(clknet_leaf_79_clk),
    .D(\sa_inst._11_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._17_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14689_ (.CLK(clknet_leaf_46_clk),
    .D(_00633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._23_ ));
 sky130_fd_sc_hd__dfxtp_1 _14690_ (.CLK(clknet_leaf_51_clk),
    .D(\sa_inst._21_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._22_ ));
 sky130_fd_sc_hd__dfxtp_1 _14691_ (.CLK(clknet_leaf_159_clk),
    .D(_00634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._02_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14692_ (.CLK(clknet_leaf_46_clk),
    .D(\sa_inst._23_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._01_ ));
 sky130_fd_sc_hd__dfxtp_4 _14693_ (.CLK(clknet_leaf_143_clk),
    .D(_00635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.WR_DATA[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14694_ (.CLK(clknet_leaf_173_clk),
    .D(\sa_inst._02_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.WR_DATA[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14695_ (.CLK(clknet_leaf_184_clk),
    .D(\sa_inst._02_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.WR_DATA[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14696_ (.CLK(clknet_leaf_161_clk),
    .D(\sa_inst._02_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.WR_DATA[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14697_ (.CLK(clknet_leaf_160_clk),
    .D(\sa_inst._02_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.WR_DATA[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14698_ (.CLK(clknet_leaf_159_clk),
    .D(\sa_inst._02_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.WR_DATA[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14699_ (.CLK(clknet_leaf_159_clk),
    .D(\sa_inst._02_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.WR_DATA[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14700_ (.CLK(clknet_leaf_159_clk),
    .D(\sa_inst._02_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.WR_DATA[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14701_ (.CLK(clknet_leaf_159_clk),
    .D(\sa_inst._02_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.WR_DATA[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14702_ (.CLK(clknet_leaf_80_clk),
    .D(_00636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sa_inst._07_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14703_ (.CLK(clknet_leaf_182_clk),
    .D(_00637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14704_ (.CLK(clknet_leaf_187_clk),
    .D(_00638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14705_ (.CLK(clknet_leaf_179_clk),
    .D(_00639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14706_ (.CLK(clknet_leaf_178_clk),
    .D(_00640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14707_ (.CLK(clknet_leaf_178_clk),
    .D(_00641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14708_ (.CLK(clknet_leaf_159_clk),
    .D(_00642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14709_ (.CLK(clknet_leaf_154_clk),
    .D(_00643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14710_ (.CLK(clknet_leaf_159_clk),
    .D(_00644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14711_ (.CLK(clknet_leaf_155_clk),
    .D(_00645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14712_ (.CLK(clknet_leaf_155_clk),
    .D(_00646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14713_ (.CLK(clknet_leaf_150_clk),
    .D(_00647_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14714_ (.CLK(clknet_leaf_149_clk),
    .D(_00648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14715_ (.CLK(clknet_leaf_148_clk),
    .D(_00649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14716_ (.CLK(clknet_leaf_147_clk),
    .D(_00650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14717_ (.CLK(clknet_leaf_148_clk),
    .D(_00651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14718_ (.CLK(clknet_leaf_4_clk),
    .D(_00652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14719_ (.CLK(clknet_leaf_4_clk),
    .D(_00653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14720_ (.CLK(clknet_leaf_4_clk),
    .D(_00654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14721_ (.CLK(clknet_leaf_6_clk),
    .D(_00655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14722_ (.CLK(clknet_leaf_1_clk),
    .D(_00656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14723_ (.CLK(clknet_leaf_190_clk),
    .D(_00657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14724_ (.CLK(clknet_leaf_190_clk),
    .D(_00658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14725_ (.CLK(clknet_leaf_188_clk),
    .D(_00659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14726_ (.CLK(clknet_leaf_189_clk),
    .D(_00660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.rMemory[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14727_ (.CLK(clknet_leaf_171_clk),
    .D(_00661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.rEmpty ));
 sky130_fd_sc_hd__dfxtp_1 _14728_ (.CLK(clknet_leaf_173_clk),
    .D(_00662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.rFull ));
 sky130_fd_sc_hd__dfxtp_4 _14729_ (.CLK(clknet_leaf_171_clk),
    .D(_00663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_1 _14730_ (.CLK(clknet_leaf_170_clk),
    .D(_00664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.rWrPtrPlus1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14731_ (.CLK(clknet_leaf_170_clk),
    .D(_00665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.rWrPtrPlus1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14732_ (.CLK(clknet_leaf_170_clk),
    .D(_00666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.rWrPtrPlus1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14733_ (.CLK(clknet_leaf_185_clk),
    .D(_00667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.rWrPtrPlus1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14734_ (.CLK(clknet_leaf_184_clk),
    .D(_00668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.rWrPtrPlus1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14735_ (.CLK(clknet_leaf_171_clk),
    .D(_00669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.WR1_ADDR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14736_ (.CLK(clknet_leaf_173_clk),
    .D(_00670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.WR1_ADDR[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14737_ (.CLK(clknet_leaf_173_clk),
    .D(_00671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.WR1_ADDR[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14738_ (.CLK(clknet_leaf_171_clk),
    .D(_00672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.WR1_ADDR[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14739_ (.CLK(clknet_leaf_171_clk),
    .D(_00673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.rWrPtr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14740_ (.CLK(clknet_leaf_183_clk),
    .D(_00674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.rRdPtrPlus1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14741_ (.CLK(clknet_leaf_183_clk),
    .D(_00675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.rRdPtrPlus1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14742_ (.CLK(clknet_leaf_183_clk),
    .D(_00676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.rRdPtrPlus1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14743_ (.CLK(clknet_leaf_184_clk),
    .D(_00677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.rRdPtrPlus1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14744_ (.CLK(clknet_leaf_184_clk),
    .D(_00678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.rRdPtrPlus1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14745_ (.CLK(clknet_leaf_171_clk),
    .D(_00679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.RD1_ADDR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14746_ (.CLK(clknet_leaf_171_clk),
    .D(_00680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.RD1_ADDR[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14747_ (.CLK(clknet_leaf_184_clk),
    .D(_00681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.RD1_ADDR[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14748_ (.CLK(clknet_leaf_184_clk),
    .D(_00682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.mem.RD1_ADDR[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14749_ (.CLK(clknet_leaf_184_clk),
    .D(_00683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fifo_inst.rRdPtr[4] ));
 sky130_fd_sc_hd__conb_1 _14750__61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net61));
 sky130_fd_sc_hd__conb_1 _14751__62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net62));
 sky130_fd_sc_hd__conb_1 _14752__63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net63));
 sky130_fd_sc_hd__conb_1 _14753__64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net64));
 sky130_fd_sc_hd__conb_1 _14754__65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net65));
 sky130_fd_sc_hd__conb_1 _14755__66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net66));
 sky130_fd_sc_hd__conb_1 _14756__67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net67));
 sky130_fd_sc_hd__conb_1 _14757__68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net68));
 sky130_fd_sc_hd__conb_1 _14758__69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net69));
 sky130_fd_sc_hd__conb_1 _14759__70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net70));
 sky130_fd_sc_hd__conb_1 _14760__71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net71));
 sky130_fd_sc_hd__conb_1 _14761__72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net72));
 sky130_fd_sc_hd__conb_1 _14762__73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net73));
 sky130_fd_sc_hd__conb_1 _14763__74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net74));
 sky130_fd_sc_hd__clkbuf_1 _14764_ (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_0_0_clk (.A(clknet_1_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_1_0_clk (.A(clknet_1_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_2_0_clk (.A(clknet_1_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_3_0_clk (.A(clknet_1_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_0_0_clk (.A(clknet_2_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_1_0_clk (.A(clknet_2_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_2_0_clk (.A(clknet_2_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_3_0_clk (.A(clknet_2_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_4_0_clk (.A(clknet_2_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_5_0_clk (.A(clknet_2_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_6_0_clk (.A(clknet_2_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_7_0_clk (.A(clknet_2_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_0_0_clk (.A(clknet_3_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_10_0_clk (.A(clknet_3_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_11_0_clk (.A(clknet_3_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_12_0_clk (.A(clknet_3_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_13_0_clk (.A(clknet_3_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_14_0_clk (.A(clknet_3_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_15_0_clk (.A(clknet_3_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_1_0_clk (.A(clknet_3_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_2_0_clk (.A(clknet_3_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_3_0_clk (.A(clknet_3_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_4_0_clk (.A(clknet_3_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_5_0_clk (.A(clknet_3_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_6_0_clk (.A(clknet_3_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_7_0_clk (.A(clknet_3_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_8_0_clk (.A(clknet_3_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_9_0_clk (.A(clknet_3_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__buf_6 input1 (.A(data_i[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input10 (.A(data_i[18]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(data_i[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(data_i[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__buf_6 input13 (.A(data_i[20]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(data_i[21]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__buf_6 input15 (.A(data_i[22]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__buf_6 input16 (.A(data_i[23]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__buf_6 input17 (.A(data_i[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(data_i[30]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(data_i[31]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(data_i[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(data_i[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(data_i[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__buf_4 input22 (.A(data_i[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__buf_6 input23 (.A(data_i[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__buf_8 input24 (.A(data_i[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(data_i[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(data_i[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__buf_4 input27 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__buf_12 input28 (.A(rtr_i),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__buf_4 input29 (.A(rts_i),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__buf_8 input3 (.A(data_i[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(data_i[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(data_i[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__buf_6 input6 (.A(data_i[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__buf_6 input7 (.A(data_i[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__buf_6 input8 (.A(data_i[16]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__buf_6 input9 (.A(data_i[17]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[0]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[10]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[11]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[12]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[13]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[14]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[15]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[16]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[17]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[18]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[19]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[1]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[20]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[21]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[22]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[23]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[2]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[3]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[4]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[5]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[6]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[7]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[8]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_o[9]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(rtr_o));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(rts_o));
 sky130_fd_sc_hd__buf_12 repeater56 (.A(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__buf_12 repeater57 (.A(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__buf_12 repeater58 (.A(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__buf_12 repeater59 (.A(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__buf_12 repeater60 (.A(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 assign data_o[24] = net61;
 assign data_o[25] = net62;
 assign data_o[26] = net63;
 assign data_o[27] = net64;
 assign data_o[28] = net65;
 assign data_o[29] = net66;
 assign data_o[30] = net67;
 assign data_o[31] = net68;
endmodule
