magic
tech sky130A
magscale 1 2
timestamp 1647539321
<< obsli1 >>
rect 1104 2159 90804 91953
<< obsm1 >>
rect 14 1980 91526 92268
<< metal2 >>
rect 3882 93328 3938 94128
rect 9034 93328 9090 94128
rect 14186 93328 14242 94128
rect 19338 93328 19394 94128
rect 24490 93328 24546 94128
rect 29642 93328 29698 94128
rect 34794 93328 34850 94128
rect 39946 93328 40002 94128
rect 45098 93328 45154 94128
rect 50250 93328 50306 94128
rect 55402 93328 55458 94128
rect 60554 93328 60610 94128
rect 65706 93328 65762 94128
rect 70858 93328 70914 94128
rect 76010 93328 76066 94128
rect 81162 93328 81218 94128
rect 86314 93328 86370 94128
rect 91466 93328 91522 94128
rect 18 0 74 800
rect 5170 0 5226 800
rect 10322 0 10378 800
rect 15474 0 15530 800
rect 20626 0 20682 800
rect 25778 0 25834 800
rect 30930 0 30986 800
rect 36082 0 36138 800
rect 41234 0 41290 800
rect 46386 0 46442 800
rect 51538 0 51594 800
rect 56690 0 56746 800
rect 61842 0 61898 800
rect 66994 0 67050 800
rect 72146 0 72202 800
rect 77298 0 77354 800
rect 82450 0 82506 800
rect 87602 0 87658 800
<< obsm2 >>
rect 20 93272 3826 93378
rect 3994 93272 8978 93378
rect 9146 93272 14130 93378
rect 14298 93272 19282 93378
rect 19450 93272 24434 93378
rect 24602 93272 29586 93378
rect 29754 93272 34738 93378
rect 34906 93272 39890 93378
rect 40058 93272 45042 93378
rect 45210 93272 50194 93378
rect 50362 93272 55346 93378
rect 55514 93272 60498 93378
rect 60666 93272 65650 93378
rect 65818 93272 70802 93378
rect 70970 93272 75954 93378
rect 76122 93272 81106 93378
rect 81274 93272 86258 93378
rect 86426 93272 91410 93378
rect 20 856 91520 93272
rect 130 800 5114 856
rect 5282 800 10266 856
rect 10434 800 15418 856
rect 15586 800 20570 856
rect 20738 800 25722 856
rect 25890 800 30874 856
rect 31042 800 36026 856
rect 36194 800 41178 856
rect 41346 800 46330 856
rect 46498 800 51482 856
rect 51650 800 56634 856
rect 56802 800 61786 856
rect 61954 800 66938 856
rect 67106 800 72090 856
rect 72258 800 77242 856
rect 77410 800 82394 856
rect 82562 800 87546 856
rect 87714 800 91520 856
<< metal3 >>
rect 0 92488 800 92608
rect 91184 88408 91984 88528
rect 0 87048 800 87168
rect 91184 82968 91984 83088
rect 0 81608 800 81728
rect 91184 77528 91984 77648
rect 0 76168 800 76288
rect 91184 72088 91984 72208
rect 0 70728 800 70848
rect 91184 66648 91984 66768
rect 0 65288 800 65408
rect 91184 61208 91984 61328
rect 0 59848 800 59968
rect 91184 55768 91984 55888
rect 0 54408 800 54528
rect 91184 50328 91984 50448
rect 0 48968 800 49088
rect 91184 44888 91984 45008
rect 0 43528 800 43648
rect 91184 39448 91984 39568
rect 0 38088 800 38208
rect 91184 34008 91984 34128
rect 0 32648 800 32768
rect 91184 28568 91984 28688
rect 0 27208 800 27328
rect 91184 23128 91984 23248
rect 0 21768 800 21888
rect 91184 17688 91984 17808
rect 0 16328 800 16448
rect 91184 12248 91984 12368
rect 0 10888 800 11008
rect 91184 6808 91984 6928
rect 0 5448 800 5568
rect 91184 1368 91984 1488
<< obsm3 >>
rect 880 92408 91184 92581
rect 800 88608 91184 92408
rect 800 88328 91104 88608
rect 800 87248 91184 88328
rect 880 86968 91184 87248
rect 800 83168 91184 86968
rect 800 82888 91104 83168
rect 800 81808 91184 82888
rect 880 81528 91184 81808
rect 800 77728 91184 81528
rect 800 77448 91104 77728
rect 800 76368 91184 77448
rect 880 76088 91184 76368
rect 800 72288 91184 76088
rect 800 72008 91104 72288
rect 800 70928 91184 72008
rect 880 70648 91184 70928
rect 800 66848 91184 70648
rect 800 66568 91104 66848
rect 800 65488 91184 66568
rect 880 65208 91184 65488
rect 800 61408 91184 65208
rect 800 61128 91104 61408
rect 800 60048 91184 61128
rect 880 59768 91184 60048
rect 800 55968 91184 59768
rect 800 55688 91104 55968
rect 800 54608 91184 55688
rect 880 54328 91184 54608
rect 800 50528 91184 54328
rect 800 50248 91104 50528
rect 800 49168 91184 50248
rect 880 48888 91184 49168
rect 800 45088 91184 48888
rect 800 44808 91104 45088
rect 800 43728 91184 44808
rect 880 43448 91184 43728
rect 800 39648 91184 43448
rect 800 39368 91104 39648
rect 800 38288 91184 39368
rect 880 38008 91184 38288
rect 800 34208 91184 38008
rect 800 33928 91104 34208
rect 800 32848 91184 33928
rect 880 32568 91184 32848
rect 800 28768 91184 32568
rect 800 28488 91104 28768
rect 800 27408 91184 28488
rect 880 27128 91184 27408
rect 800 23328 91184 27128
rect 800 23048 91104 23328
rect 800 21968 91184 23048
rect 880 21688 91184 21968
rect 800 17888 91184 21688
rect 800 17608 91104 17888
rect 800 16528 91184 17608
rect 880 16248 91184 16528
rect 800 12448 91184 16248
rect 800 12168 91104 12448
rect 800 11088 91184 12168
rect 880 10808 91184 11088
rect 800 7008 91184 10808
rect 800 6728 91104 7008
rect 800 5648 91184 6728
rect 880 5368 91184 5648
rect 800 1568 91184 5368
rect 800 1395 91104 1568
<< metal4 >>
rect 4208 2128 4528 91984
rect 19568 2128 19888 91984
rect 34928 2128 35248 91984
rect 50288 2128 50608 91984
rect 65648 2128 65968 91984
rect 81008 2128 81328 91984
<< obsm4 >>
rect 14227 2347 19488 88365
rect 19968 2347 34848 88365
rect 35328 2347 50208 88365
rect 50688 2347 65568 88365
rect 66048 2347 80928 88365
rect 81408 2347 86421 88365
<< metal5 >>
rect 1104 81888 90804 82208
rect 1104 66570 90804 66890
rect 1104 51252 90804 51572
rect 1104 35934 90804 36254
rect 1104 20616 90804 20936
rect 1104 5298 90804 5618
<< labels >>
rlabel metal5 s 1104 20616 90804 20936 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 51252 90804 51572 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 81888 90804 82208 6 VGND
port 1 nsew ground input
rlabel metal4 s 19568 2128 19888 91984 6 VGND
port 1 nsew ground input
rlabel metal4 s 50288 2128 50608 91984 6 VGND
port 1 nsew ground input
rlabel metal4 s 81008 2128 81328 91984 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 5298 90804 5618 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 35934 90804 36254 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 66570 90804 66890 6 VPWR
port 2 nsew power input
rlabel metal4 s 4208 2128 4528 91984 6 VPWR
port 2 nsew power input
rlabel metal4 s 34928 2128 35248 91984 6 VPWR
port 2 nsew power input
rlabel metal4 s 65648 2128 65968 91984 6 VPWR
port 2 nsew power input
rlabel metal2 s 20626 0 20682 800 6 clk
port 3 nsew signal input
rlabel metal3 s 91184 39448 91984 39568 6 data_i[0]
port 4 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 data_i[10]
port 5 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 data_i[11]
port 6 nsew signal input
rlabel metal2 s 9034 93328 9090 94128 6 data_i[12]
port 7 nsew signal input
rlabel metal3 s 91184 61208 91984 61328 6 data_i[13]
port 8 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 data_i[14]
port 9 nsew signal input
rlabel metal3 s 91184 12248 91984 12368 6 data_i[15]
port 10 nsew signal input
rlabel metal3 s 91184 17688 91984 17808 6 data_i[16]
port 11 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 data_i[17]
port 12 nsew signal input
rlabel metal3 s 91184 72088 91984 72208 6 data_i[18]
port 13 nsew signal input
rlabel metal3 s 0 92488 800 92608 6 data_i[19]
port 14 nsew signal input
rlabel metal3 s 91184 66648 91984 66768 6 data_i[1]
port 15 nsew signal input
rlabel metal3 s 91184 6808 91984 6928 6 data_i[20]
port 16 nsew signal input
rlabel metal2 s 29642 93328 29698 94128 6 data_i[21]
port 17 nsew signal input
rlabel metal3 s 91184 28568 91984 28688 6 data_i[22]
port 18 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 data_i[23]
port 19 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 data_i[24]
port 20 nsew signal input
rlabel metal3 s 91184 55768 91984 55888 6 data_i[25]
port 21 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 data_i[26]
port 22 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 data_i[27]
port 23 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 data_i[28]
port 24 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 data_i[29]
port 25 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 data_i[2]
port 26 nsew signal input
rlabel metal2 s 39946 93328 40002 94128 6 data_i[30]
port 27 nsew signal input
rlabel metal2 s 70858 93328 70914 94128 6 data_i[31]
port 28 nsew signal input
rlabel metal2 s 19338 93328 19394 94128 6 data_i[3]
port 29 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 data_i[4]
port 30 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 data_i[5]
port 31 nsew signal input
rlabel metal2 s 91466 93328 91522 94128 6 data_i[6]
port 32 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 data_i[7]
port 33 nsew signal input
rlabel metal2 s 50250 93328 50306 94128 6 data_i[8]
port 34 nsew signal input
rlabel metal3 s 91184 88408 91984 88528 6 data_i[9]
port 35 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 data_o[0]
port 36 nsew signal output
rlabel metal2 s 45098 93328 45154 94128 6 data_o[10]
port 37 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 data_o[11]
port 38 nsew signal output
rlabel metal3 s 91184 23128 91984 23248 6 data_o[12]
port 39 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 data_o[13]
port 40 nsew signal output
rlabel metal3 s 91184 34008 91984 34128 6 data_o[14]
port 41 nsew signal output
rlabel metal2 s 60554 93328 60610 94128 6 data_o[15]
port 42 nsew signal output
rlabel metal2 s 65706 93328 65762 94128 6 data_o[16]
port 43 nsew signal output
rlabel metal2 s 3882 93328 3938 94128 6 data_o[17]
port 44 nsew signal output
rlabel metal2 s 18 0 74 800 6 data_o[18]
port 45 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 data_o[19]
port 46 nsew signal output
rlabel metal2 s 55402 93328 55458 94128 6 data_o[1]
port 47 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 data_o[20]
port 48 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 data_o[21]
port 49 nsew signal output
rlabel metal2 s 34794 93328 34850 94128 6 data_o[22]
port 50 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 data_o[23]
port 51 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 data_o[24]
port 52 nsew signal output
rlabel metal3 s 91184 82968 91984 83088 6 data_o[25]
port 53 nsew signal output
rlabel metal2 s 86314 93328 86370 94128 6 data_o[26]
port 54 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 data_o[27]
port 55 nsew signal output
rlabel metal3 s 91184 77528 91984 77648 6 data_o[28]
port 56 nsew signal output
rlabel metal3 s 91184 1368 91984 1488 6 data_o[29]
port 57 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 data_o[2]
port 58 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 data_o[30]
port 59 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 data_o[31]
port 60 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 data_o[3]
port 61 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 data_o[4]
port 62 nsew signal output
rlabel metal3 s 91184 50328 91984 50448 6 data_o[5]
port 63 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 data_o[6]
port 64 nsew signal output
rlabel metal2 s 81162 93328 81218 94128 6 data_o[7]
port 65 nsew signal output
rlabel metal2 s 76010 93328 76066 94128 6 data_o[8]
port 66 nsew signal output
rlabel metal2 s 14186 93328 14242 94128 6 data_o[9]
port 67 nsew signal output
rlabel metal2 s 24490 93328 24546 94128 6 rst_n
port 68 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 rtr_i
port 69 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 rtr_o
port 70 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 rts_i
port 71 nsew signal input
rlabel metal3 s 91184 44888 91984 45008 6 rts_o
port 72 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 91984 94128
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 23504280
string GDS_FILE /openlane/designs/teras/runs/RUN_2022.03.17_17.43.33/results/finishing/teras.magic.gds
string GDS_START 1108954
<< end >>

